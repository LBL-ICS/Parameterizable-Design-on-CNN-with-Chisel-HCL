module full_subber(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s,
  output       io_out_c
);
  wire [8:0] _result_T = io_in_a - io_in_b; // @[Arithmetic.scala 70:23]
  wire [9:0] _result_T_2 = _result_T - 9'h0; // @[Arithmetic.scala 70:34]
  wire [8:0] result = _result_T_2[8:0]; // @[Arithmetic.scala 69:22 70:12]
  assign io_out_s = result[7:0]; // @[Arithmetic.scala 71:23]
  assign io_out_c = result[8]; // @[Arithmetic.scala 72:23]
endmodule
module twoscomplement(
  input  [7:0] io_in,
  output [7:0] io_out
);
  wire [7:0] x = ~io_in; // @[Arithmetic.scala 26:10]
  assign io_out = x + 8'h1; // @[Arithmetic.scala 27:17]
endmodule
module full_adder(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [23:0] io_out_s,
  output        io_out_c
);
  wire [24:0] _result_T = io_in_a + io_in_b; // @[Arithmetic.scala 56:23]
  wire [25:0] _result_T_1 = {{1'd0}, _result_T}; // @[Arithmetic.scala 56:34]
  wire [24:0] result = _result_T_1[24:0]; // @[Arithmetic.scala 55:22 56:12]
  assign io_out_s = result[23:0]; // @[Arithmetic.scala 57:23]
  assign io_out_c = result[24]; // @[Arithmetic.scala 58:23]
endmodule
module twoscomplement_1(
  input  [23:0] io_in,
  output [23:0] io_out
);
  wire [23:0] x = ~io_in; // @[Arithmetic.scala 26:10]
  assign io_out = x + 24'h1; // @[Arithmetic.scala 27:17]
endmodule
module shifter(
  input  [23:0] io_in_a,
  input  [4:0]  io_in_b,
  output [23:0] io_out_s
);
  wire [23:0] _result_T = io_in_a >> io_in_b; // @[Arithmetic.scala 40:25]
  wire [54:0] _GEN_0 = {{31'd0}, _result_T}; // @[Arithmetic.scala 39:26 40:14 42:14]
  assign io_out_s = _GEN_0[23:0]; // @[Arithmetic.scala 37:22]
endmodule
module leadingOneDetector(
  input  [23:0] io_in,
  output [4:0]  io_out
);
  wire [1:0] _hotValue_T = io_in[1] ? 2'h2 : 2'h1; // @[Mux.scala 47:70]
  wire [1:0] _hotValue_T_1 = io_in[2] ? 2'h3 : _hotValue_T; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_2 = io_in[3] ? 3'h4 : {{1'd0}, _hotValue_T_1}; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_3 = io_in[4] ? 3'h5 : _hotValue_T_2; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_4 = io_in[5] ? 3'h6 : _hotValue_T_3; // @[Mux.scala 47:70]
  wire [2:0] _hotValue_T_5 = io_in[6] ? 3'h7 : _hotValue_T_4; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_6 = io_in[7] ? 4'h8 : {{1'd0}, _hotValue_T_5}; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_7 = io_in[8] ? 4'h9 : _hotValue_T_6; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_8 = io_in[9] ? 4'ha : _hotValue_T_7; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_9 = io_in[10] ? 4'hb : _hotValue_T_8; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_10 = io_in[11] ? 4'hc : _hotValue_T_9; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_11 = io_in[12] ? 4'hd : _hotValue_T_10; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_12 = io_in[13] ? 4'he : _hotValue_T_11; // @[Mux.scala 47:70]
  wire [3:0] _hotValue_T_13 = io_in[14] ? 4'hf : _hotValue_T_12; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_14 = io_in[15] ? 5'h10 : {{1'd0}, _hotValue_T_13}; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_15 = io_in[16] ? 5'h11 : _hotValue_T_14; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_16 = io_in[17] ? 5'h12 : _hotValue_T_15; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_17 = io_in[18] ? 5'h13 : _hotValue_T_16; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_18 = io_in[19] ? 5'h14 : _hotValue_T_17; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_19 = io_in[20] ? 5'h15 : _hotValue_T_18; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_20 = io_in[21] ? 5'h16 : _hotValue_T_19; // @[Mux.scala 47:70]
  wire [4:0] _hotValue_T_21 = io_in[22] ? 5'h17 : _hotValue_T_20; // @[Mux.scala 47:70]
  assign io_out = io_in[23] ? 5'h18 : _hotValue_T_21; // @[Mux.scala 47:70]
endmodule
module FP_adder(
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
  wire [7:0] subber_io_in_a; // @[FPArithmetic.scala 72:24]
  wire [7:0] subber_io_in_b; // @[FPArithmetic.scala 72:24]
  wire [7:0] subber_io_out_s; // @[FPArithmetic.scala 72:24]
  wire  subber_io_out_c; // @[FPArithmetic.scala 72:24]
  wire [7:0] complement_io_in; // @[FPArithmetic.scala 78:28]
  wire [7:0] complement_io_out; // @[FPArithmetic.scala 78:28]
  wire [23:0] adder_io_in_a; // @[FPArithmetic.scala 82:23]
  wire [23:0] adder_io_in_b; // @[FPArithmetic.scala 82:23]
  wire [23:0] adder_io_out_s; // @[FPArithmetic.scala 82:23]
  wire  adder_io_out_c; // @[FPArithmetic.scala 82:23]
  wire [23:0] complementN_0_io_in; // @[FPArithmetic.scala 88:31]
  wire [23:0] complementN_0_io_out; // @[FPArithmetic.scala 88:31]
  wire [23:0] complementN_1_io_in; // @[FPArithmetic.scala 90:31]
  wire [23:0] complementN_1_io_out; // @[FPArithmetic.scala 90:31]
  wire [23:0] shifter_io_in_a; // @[FPArithmetic.scala 94:25]
  wire [4:0] shifter_io_in_b; // @[FPArithmetic.scala 94:25]
  wire [23:0] shifter_io_out_s; // @[FPArithmetic.scala 94:25]
  wire [23:0] complementN_2_io_in; // @[FPArithmetic.scala 139:31]
  wire [23:0] complementN_2_io_out; // @[FPArithmetic.scala 139:31]
  wire [23:0] leadingOneFinder_io_in; // @[FPArithmetic.scala 159:34]
  wire [4:0] leadingOneFinder_io_out; // @[FPArithmetic.scala 159:34]
  wire [7:0] subber2_io_in_a; // @[FPArithmetic.scala 161:25]
  wire [7:0] subber2_io_in_b; // @[FPArithmetic.scala 161:25]
  wire [7:0] subber2_io_out_s; // @[FPArithmetic.scala 161:25]
  wire  subber2_io_out_c; // @[FPArithmetic.scala 161:25]
  wire  sign_0 = io_in_a[31]; // @[FPArithmetic.scala 34:23]
  wire  sign_1 = io_in_b[31]; // @[FPArithmetic.scala 35:23]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FPArithmetic.scala 39:62]
  wire [8:0] _GEN_31 = {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 39:34]
  wire [8:0] _GEN_0 = _GEN_31 > _T_2 ? _T_2 : {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 39:68 40:14 42:14]
  wire [8:0] _GEN_32 = {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 44:34]
  wire [8:0] _GEN_1 = _GEN_32 > _T_2 ? _T_2 : {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 44:68 45:14 47:14]
  wire [22:0] frac_0 = io_in_a[22:0]; // @[FPArithmetic.scala 52:23]
  wire [22:0] frac_1 = io_in_b[22:0]; // @[FPArithmetic.scala 53:23]
  wire [23:0] whole_frac_0 = {1'h1,frac_0}; // @[FPArithmetic.scala 57:26]
  wire [23:0] whole_frac_1 = {1'h1,frac_1}; // @[FPArithmetic.scala 58:26]
  wire [7:0] exp_1 = _GEN_1[7:0]; // @[FPArithmetic.scala 38:19]
  wire [7:0] exp_0 = _GEN_0[7:0]; // @[FPArithmetic.scala 38:19]
  wire [7:0] out_exp = subber_io_out_c ? exp_1 : exp_0; // @[FPArithmetic.scala 100:34 101:15 111:15]
  wire [7:0] sub_exp = subber_io_out_c ? complement_io_out : subber_io_out_s; // @[FPArithmetic.scala 100:34 102:15 112:15]
  wire  out_s = subber_io_out_c ? sign_1 : sign_0; // @[FPArithmetic.scala 100:34 103:13 113:13]
  wire [22:0] out_frac = subber_io_out_c ? frac_1 : frac_0; // @[FPArithmetic.scala 100:34 104:16 114:16]
  wire [23:0] _GEN_8 = subber_io_out_c ? shifter_io_out_s : whole_frac_0; // @[FPArithmetic.scala 100:34 108:21 83:19]
  wire [23:0] _GEN_9 = subber_io_out_c ? whole_frac_1 : shifter_io_out_s; // @[FPArithmetic.scala 100:34 84:19 118:21]
  wire  _new_s_T = ~adder_io_out_c; // @[FPArithmetic.scala 134:15]
  wire  _D_T_1 = sign_0 ^ sign_1; // @[FPArithmetic.scala 147:39]
  wire  D = _new_s_T | sign_0 ^ sign_1; // @[FPArithmetic.scala 147:28]
  wire  E = _new_s_T & ~adder_io_out_s[23] | _new_s_T & ~_D_T_1 | adder_io_out_c & adder_io_out_s[23] & _D_T_1; // @[FPArithmetic.scala 150:99]
  wire  _GEN_25 = sub_exp >= 8'h17 ? out_s : ~adder_io_out_c & sign_0 | sign_0 & sign_1 | ~adder_io_out_c & sign_1; // @[FPArithmetic.scala 134:11 166:33 167:13]
  wire  new_s = io_in_a[30:0] == 31'h0 & io_in_b[30:0] == 31'h0 ? 1'h0 : _GEN_25; // @[FPArithmetic.scala 194:62 195:13]
  wire [23:0] adder_result = new_s & sign_0 != sign_1 ? complementN_2_io_out : adder_io_out_s; // @[FPArithmetic.scala 153:18 154:47 155:20]
  wire [4:0] _subber2_io_in_b_T_1 = 5'h18 - leadingOneFinder_io_out; // @[FPArithmetic.scala 163:42]
  wire [8:0] _GEN_33 = {{1'd0}, out_exp}; // @[FPArithmetic.scala 174:20]
  wire [23:0] _new_out_frac_T_2 = 24'h800000 - 24'h1; // @[FPArithmetic.scala 176:51]
  wire [7:0] _new_out_exp_T_3 = out_exp + 8'h1; // @[FPArithmetic.scala 178:32]
  wire [8:0] _GEN_13 = _GEN_33 == _T_2 ? _T_2 : {{1'd0}, _new_out_exp_T_3}; // @[FPArithmetic.scala 174:56 175:21 178:21]
  wire [23:0] _GEN_14 = _GEN_33 == _T_2 ? _new_out_frac_T_2 : {{1'd0}, adder_result[23:1]}; // @[FPArithmetic.scala 174:56 176:22 179:22]
  wire [53:0] _GEN_2 = {{31'd0}, adder_result[22:0]}; // @[FPArithmetic.scala 190:57]
  wire [53:0] _new_out_frac_T_7 = _GEN_2 << _subber2_io_in_b_T_1; // @[FPArithmetic.scala 190:57]
  wire [7:0] _GEN_15 = subber2_io_out_c ? 8'h1 : subber2_io_out_s; // @[FPArithmetic.scala 185:39 186:23 189:23]
  wire [53:0] _GEN_16 = subber2_io_out_c ? 54'h0 : _new_out_frac_T_7; // @[FPArithmetic.scala 185:39 187:24 190:24]
  wire [7:0] _GEN_17 = leadingOneFinder_io_out == 5'h1 & adder_result == 24'h0 & (_D_T_1 & io_in_a[30:0] == io_in_b[30:0
    ]) ? 8'h0 : _GEN_15; // @[FPArithmetic.scala 182:141 183:21]
  wire [53:0] _GEN_18 = leadingOneFinder_io_out == 5'h1 & adder_result == 24'h0 & (_D_T_1 & io_in_a[30:0] == io_in_b[30:
    0]) ? 54'h0 : _GEN_16; // @[FPArithmetic.scala 182:141 135:18]
  wire [7:0] _GEN_19 = D ? _GEN_17 : 8'h0; // @[FPArithmetic.scala 136:17 181:26]
  wire [53:0] _GEN_20 = D ? _GEN_18 : 54'h0; // @[FPArithmetic.scala 135:18 181:26]
  wire [8:0] _GEN_21 = ~D ? _GEN_13 : {{1'd0}, _GEN_19}; // @[FPArithmetic.scala 173:26]
  wire [53:0] _GEN_22 = ~D ? {{30'd0}, _GEN_14} : _GEN_20; // @[FPArithmetic.scala 173:26]
  wire [8:0] _GEN_23 = E ? {{1'd0}, out_exp} : _GEN_21; // @[FPArithmetic.scala 170:26 171:19]
  wire [53:0] _GEN_24 = E ? {{31'd0}, adder_result[22:0]} : _GEN_22; // @[FPArithmetic.scala 170:26 172:20]
  wire [53:0] _GEN_26 = sub_exp >= 8'h17 ? {{31'd0}, out_frac} : _GEN_24; // @[FPArithmetic.scala 166:33 168:20]
  wire [8:0] _GEN_27 = sub_exp >= 8'h17 ? {{1'd0}, out_exp} : _GEN_23; // @[FPArithmetic.scala 166:33 169:19]
  wire [8:0] _GEN_29 = io_in_a[30:0] == 31'h0 & io_in_b[30:0] == 31'h0 ? 9'h0 : _GEN_27; // @[FPArithmetic.scala 194:62 196:19]
  wire [53:0] _GEN_30 = io_in_a[30:0] == 31'h0 & io_in_b[30:0] == 31'h0 ? 54'h0 : _GEN_26; // @[FPArithmetic.scala 194:62 197:20]
  wire [7:0] new_out_exp = _GEN_29[7:0]; // @[FPArithmetic.scala 133:27]
  wire [8:0] _io_out_s_T = {new_s,new_out_exp}; // @[FPArithmetic.scala 201:23]
  wire [22:0] new_out_frac = _GEN_30[22:0]; // @[FPArithmetic.scala 132:28]
  full_subber subber ( // @[FPArithmetic.scala 72:24]
    .io_in_a(subber_io_in_a),
    .io_in_b(subber_io_in_b),
    .io_out_s(subber_io_out_s),
    .io_out_c(subber_io_out_c)
  );
  twoscomplement complement ( // @[FPArithmetic.scala 78:28]
    .io_in(complement_io_in),
    .io_out(complement_io_out)
  );
  full_adder adder ( // @[FPArithmetic.scala 82:23]
    .io_in_a(adder_io_in_a),
    .io_in_b(adder_io_in_b),
    .io_out_s(adder_io_out_s),
    .io_out_c(adder_io_out_c)
  );
  twoscomplement_1 complementN_0 ( // @[FPArithmetic.scala 88:31]
    .io_in(complementN_0_io_in),
    .io_out(complementN_0_io_out)
  );
  twoscomplement_1 complementN_1 ( // @[FPArithmetic.scala 90:31]
    .io_in(complementN_1_io_in),
    .io_out(complementN_1_io_out)
  );
  shifter shifter ( // @[FPArithmetic.scala 94:25]
    .io_in_a(shifter_io_in_a),
    .io_in_b(shifter_io_in_b),
    .io_out_s(shifter_io_out_s)
  );
  twoscomplement_1 complementN_2 ( // @[FPArithmetic.scala 139:31]
    .io_in(complementN_2_io_in),
    .io_out(complementN_2_io_out)
  );
  leadingOneDetector leadingOneFinder ( // @[FPArithmetic.scala 159:34]
    .io_in(leadingOneFinder_io_in),
    .io_out(leadingOneFinder_io_out)
  );
  full_subber subber2 ( // @[FPArithmetic.scala 161:25]
    .io_in_a(subber2_io_in_a),
    .io_in_b(subber2_io_in_b),
    .io_out_s(subber2_io_out_s),
    .io_out_c(subber2_io_out_c)
  );
  assign io_out_s = {_io_out_s_T,new_out_frac}; // @[FPArithmetic.scala 201:38]
  assign subber_io_in_a = _GEN_0[7:0]; // @[FPArithmetic.scala 38:19]
  assign subber_io_in_b = _GEN_1[7:0]; // @[FPArithmetic.scala 38:19]
  assign complement_io_in = subber_io_out_s; // @[FPArithmetic.scala 79:22]
  assign adder_io_in_a = sign_0 & ~sign_1 ? complementN_0_io_out : _GEN_8; // @[FPArithmetic.scala 123:45 124:21]
  assign adder_io_in_b = sign_1 & ~sign_0 ? complementN_1_io_out : _GEN_9; // @[FPArithmetic.scala 127:45 128:21]
  assign complementN_0_io_in = subber_io_out_c ? shifter_io_out_s : whole_frac_0; // @[FPArithmetic.scala 100:34 108:21 83:19]
  assign complementN_1_io_in = subber_io_out_c ? whole_frac_1 : shifter_io_out_s; // @[FPArithmetic.scala 100:34 84:19 118:21]
  assign shifter_io_in_a = subber_io_out_c ? whole_frac_0 : whole_frac_1; // @[FPArithmetic.scala 100:34 105:23 115:23]
  assign shifter_io_in_b = sub_exp[4:0];
  assign complementN_2_io_in = adder_io_out_s; // @[FPArithmetic.scala 140:25]
  assign leadingOneFinder_io_in = new_s & sign_0 != sign_1 ? complementN_2_io_out : adder_io_out_s; // @[FPArithmetic.scala 153:18 154:47 155:20]
  assign subber2_io_in_a = subber_io_out_c ? exp_1 : exp_0; // @[FPArithmetic.scala 100:34 101:15 111:15]
  assign subber2_io_in_b = {{3'd0}, _subber2_io_in_b_T_1}; // @[FPArithmetic.scala 163:21]
endmodule
module multiplier(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [47:0] io_out_s
);
  assign io_out_s = io_in_a * io_in_b; // @[Arithmetic.scala 82:23]
endmodule
module full_adder_1(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s
);
  wire [8:0] _result_T = io_in_a + io_in_b; // @[Arithmetic.scala 56:23]
  wire [9:0] _result_T_1 = {{1'd0}, _result_T}; // @[Arithmetic.scala 56:34]
  wire [8:0] result = _result_T_1[8:0]; // @[Arithmetic.scala 55:22 56:12]
  assign io_out_s = result[7:0]; // @[Arithmetic.scala 57:23]
endmodule
module FP_multiplier(
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
  wire [23:0] multiplier_io_in_a; // @[FPArithmetic.scala 283:28]
  wire [23:0] multiplier_io_in_b; // @[FPArithmetic.scala 283:28]
  wire [47:0] multiplier_io_out_s; // @[FPArithmetic.scala 283:28]
  wire [7:0] subber_io_in_a; // @[FPArithmetic.scala 288:24]
  wire [7:0] subber_io_in_b; // @[FPArithmetic.scala 288:24]
  wire [7:0] subber_io_out_s; // @[FPArithmetic.scala 288:24]
  wire  subber_io_out_c; // @[FPArithmetic.scala 288:24]
  wire [7:0] complementN_io_in; // @[FPArithmetic.scala 294:29]
  wire [7:0] complementN_io_out; // @[FPArithmetic.scala 294:29]
  wire [7:0] adderN_io_in_a; // @[FPArithmetic.scala 298:24]
  wire [7:0] adderN_io_in_b; // @[FPArithmetic.scala 298:24]
  wire [7:0] adderN_io_out_s; // @[FPArithmetic.scala 298:24]
  wire  s_0 = io_in_a[31]; // @[FPArithmetic.scala 248:20]
  wire  s_1 = io_in_b[31]; // @[FPArithmetic.scala 249:20]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FPArithmetic.scala 253:62]
  wire [8:0] _GEN_11 = {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 253:34]
  wire [8:0] _GEN_0 = _GEN_11 > _T_2 ? _T_2 : {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 253:68 254:14 256:14]
  wire [8:0] _GEN_12 = {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 258:34]
  wire [8:0] _GEN_1 = _GEN_12 > _T_2 ? _T_2 : {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 258:68 259:14 261:14]
  wire [22:0] exp_check_0 = {{15'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 264:25 265:18]
  wire [22:0] _cond_holder_T_1 = exp_check_0 + 23'h1; // @[FPArithmetic.scala 269:34]
  wire [22:0] exp_check_1 = {{15'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 264:25 266:18]
  wire [22:0] _cond_holder_T_3 = 23'h7f - exp_check_1; // @[FPArithmetic.scala 269:80]
  wire [22:0] _cond_holder_T_4 = ~_cond_holder_T_3; // @[FPArithmetic.scala 269:42]
  wire [22:0] _cond_holder_T_6 = _cond_holder_T_1 + _cond_holder_T_4; // @[FPArithmetic.scala 269:40]
  wire [22:0] frac_0 = io_in_a[22:0]; // @[FPArithmetic.scala 273:23]
  wire [22:0] frac_1 = io_in_b[22:0]; // @[FPArithmetic.scala 274:23]
  wire  new_s = s_0 ^ s_1; // @[FPArithmetic.scala 305:19]
  wire [7:0] _new_exp_T_1 = adderN_io_out_s + 8'h1; // @[FPArithmetic.scala 316:34]
  wire [22:0] _cond_holder_T_8 = exp_check_0 + 23'h2; // @[FPArithmetic.scala 318:36]
  wire [22:0] _cond_holder_T_13 = _cond_holder_T_8 + _cond_holder_T_4; // @[FPArithmetic.scala 318:42]
  wire [23:0] _new_mant_T_2 = {multiplier_io_out_s[46:24], 1'h0}; // @[FPArithmetic.scala 324:73]
  wire [7:0] _GEN_2 = multiplier_io_out_s[47] ? _new_exp_T_1 : adderN_io_out_s; // @[FPArithmetic.scala 315:60 316:15 321:15]
  wire [22:0] cond_holder = multiplier_io_out_s[47] ? _cond_holder_T_13 : _cond_holder_T_6; // @[FPArithmetic.scala 315:60 318:19 323:19]
  wire [23:0] _GEN_5 = multiplier_io_out_s[47] ? {{1'd0}, multiplier_io_out_s[46:24]} : _new_mant_T_2; // @[FPArithmetic.scala 315:60 319:16 324:16]
  wire [22:0] _T_12 = ~cond_holder; // @[FPArithmetic.scala 327:51]
  wire [22:0] _T_14 = 23'h1 + _T_12; // @[FPArithmetic.scala 327:49]
  wire [22:0] _GEN_13 = {{14'd0}, _T_2}; // @[FPArithmetic.scala 327:42]
  wire [8:0] _GEN_6 = cond_holder > _GEN_13 ? _T_2 : {{1'd0}, _GEN_2}; // @[FPArithmetic.scala 332:63 333:17]
  wire [8:0] _GEN_8 = _GEN_13 >= _T_14 ? 9'h1 : _GEN_6; // @[FPArithmetic.scala 327:67 328:15]
  wire [7:0] new_exp = _GEN_8[7:0]; // @[FPArithmetic.scala 308:23]
  wire [23:0] _new_mant_T_4 = 24'h800000 - 24'h1; // @[FPArithmetic.scala 334:47]
  wire [23:0] _GEN_7 = cond_holder > _GEN_13 ? _new_mant_T_4 : _GEN_5; // @[FPArithmetic.scala 332:63 334:18]
  wire [23:0] _GEN_9 = _GEN_13 >= _T_14 ? 24'h0 : _GEN_7; // @[FPArithmetic.scala 327:67 329:16]
  wire [22:0] new_mant = _GEN_9[22:0]; // @[FPArithmetic.scala 310:24]
  wire [31:0] _io_out_s_T_1 = {new_s,new_exp,new_mant}; // @[FPArithmetic.scala 330:36]
  wire [7:0] exp_0 = _GEN_0[7:0]; // @[FPArithmetic.scala 252:19]
  wire [7:0] exp_1 = _GEN_1[7:0]; // @[FPArithmetic.scala 252:19]
  multiplier multiplier ( // @[FPArithmetic.scala 283:28]
    .io_in_a(multiplier_io_in_a),
    .io_in_b(multiplier_io_in_b),
    .io_out_s(multiplier_io_out_s)
  );
  full_subber subber ( // @[FPArithmetic.scala 288:24]
    .io_in_a(subber_io_in_a),
    .io_in_b(subber_io_in_b),
    .io_out_s(subber_io_out_s),
    .io_out_c(subber_io_out_c)
  );
  twoscomplement complementN ( // @[FPArithmetic.scala 294:29]
    .io_in(complementN_io_in),
    .io_out(complementN_io_out)
  );
  full_adder_1 adderN ( // @[FPArithmetic.scala 298:24]
    .io_in_a(adderN_io_in_a),
    .io_in_b(adderN_io_in_b),
    .io_out_s(adderN_io_out_s)
  );
  assign io_out_s = exp_0 == 8'h0 | exp_1 == 8'h0 ? 32'h0 : _io_out_s_T_1; // @[FPArithmetic.scala 337:43 338:16 340:16]
  assign multiplier_io_in_a = {1'h1,frac_0}; // @[FPArithmetic.scala 278:24]
  assign multiplier_io_in_b = {1'h1,frac_1}; // @[FPArithmetic.scala 279:24]
  assign subber_io_in_a = 8'h7f; // @[FPArithmetic.scala 289:20]
  assign subber_io_in_b = _GEN_1[7:0]; // @[FPArithmetic.scala 252:19]
  assign complementN_io_in = subber_io_out_s; // @[FPArithmetic.scala 295:23]
  assign adderN_io_in_a = _GEN_0[7:0]; // @[FPArithmetic.scala 252:19]
  assign adderN_io_in_b = complementN_io_out; // @[FPArithmetic.scala 300:20]
endmodule
module FP_multiply_sum(
  input  [31:0] io_in_a_0,
  input  [31:0] io_in_a_1,
  input  [31:0] io_in_a_2,
  input  [31:0] io_in_a_3,
  input  [31:0] io_in_a_4,
  input  [31:0] io_in_a_5,
  input  [31:0] io_in_a_6,
  input  [31:0] io_in_a_7,
  input  [31:0] io_in_a_8,
  output [31:0] io_out_s
);
  wire [31:0] FP_multipliers_0_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_0_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_0_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_1_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_1_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_1_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_2_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_2_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_2_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_3_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_3_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_3_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_4_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_4_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_4_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_5_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_5_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_5_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_6_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_6_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_6_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_7_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_7_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_7_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_8_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_8_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_8_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_adders_0_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_0_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_0_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_1_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_1_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_1_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_2_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_2_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_2_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_3_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_3_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_3_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_4_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_4_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_4_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_5_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_5_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_5_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_6_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_6_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_6_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_7_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_7_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_7_io_out_s; // @[FPArithmetic.scala 630:28]
  FP_multiplier FP_multipliers_0 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_0_io_in_a),
    .io_in_b(FP_multipliers_0_io_in_b),
    .io_out_s(FP_multipliers_0_io_out_s)
  );
  FP_multiplier FP_multipliers_1 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_1_io_in_a),
    .io_in_b(FP_multipliers_1_io_in_b),
    .io_out_s(FP_multipliers_1_io_out_s)
  );
  FP_multiplier FP_multipliers_2 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_2_io_in_a),
    .io_in_b(FP_multipliers_2_io_in_b),
    .io_out_s(FP_multipliers_2_io_out_s)
  );
  FP_multiplier FP_multipliers_3 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_3_io_in_a),
    .io_in_b(FP_multipliers_3_io_in_b),
    .io_out_s(FP_multipliers_3_io_out_s)
  );
  FP_multiplier FP_multipliers_4 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_4_io_in_a),
    .io_in_b(FP_multipliers_4_io_in_b),
    .io_out_s(FP_multipliers_4_io_out_s)
  );
  FP_multiplier FP_multipliers_5 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_5_io_in_a),
    .io_in_b(FP_multipliers_5_io_in_b),
    .io_out_s(FP_multipliers_5_io_out_s)
  );
  FP_multiplier FP_multipliers_6 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_6_io_in_a),
    .io_in_b(FP_multipliers_6_io_in_b),
    .io_out_s(FP_multipliers_6_io_out_s)
  );
  FP_multiplier FP_multipliers_7 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_7_io_in_a),
    .io_in_b(FP_multipliers_7_io_in_b),
    .io_out_s(FP_multipliers_7_io_out_s)
  );
  FP_multiplier FP_multipliers_8 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_8_io_in_a),
    .io_in_b(FP_multipliers_8_io_in_b),
    .io_out_s(FP_multipliers_8_io_out_s)
  );
  FP_adder FP_adders_0 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_0_io_in_a),
    .io_in_b(FP_adders_0_io_in_b),
    .io_out_s(FP_adders_0_io_out_s)
  );
  FP_adder FP_adders_1 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_1_io_in_a),
    .io_in_b(FP_adders_1_io_in_b),
    .io_out_s(FP_adders_1_io_out_s)
  );
  FP_adder FP_adders_2 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_2_io_in_a),
    .io_in_b(FP_adders_2_io_in_b),
    .io_out_s(FP_adders_2_io_out_s)
  );
  FP_adder FP_adders_3 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_3_io_in_a),
    .io_in_b(FP_adders_3_io_in_b),
    .io_out_s(FP_adders_3_io_out_s)
  );
  FP_adder FP_adders_4 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_4_io_in_a),
    .io_in_b(FP_adders_4_io_in_b),
    .io_out_s(FP_adders_4_io_out_s)
  );
  FP_adder FP_adders_5 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_5_io_in_a),
    .io_in_b(FP_adders_5_io_in_b),
    .io_out_s(FP_adders_5_io_out_s)
  );
  FP_adder FP_adders_6 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_6_io_in_a),
    .io_in_b(FP_adders_6_io_in_b),
    .io_out_s(FP_adders_6_io_out_s)
  );
  FP_adder FP_adders_7 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_7_io_in_a),
    .io_in_b(FP_adders_7_io_in_b),
    .io_out_s(FP_adders_7_io_out_s)
  );
  assign io_out_s = FP_adders_7_io_out_s; // @[FPArithmetic.scala 693:14]
  assign FP_multipliers_0_io_in_a = io_in_a_0; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_0_io_in_b = 32'h3db81d70; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_1_io_in_a = io_in_a_1; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_1_io_in_b = 32'h3ff49518; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_2_io_in_a = io_in_a_2; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_2_io_in_b = 32'h3e7ae140; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_3_io_in_a = io_in_a_3; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_3_io_in_b = 32'h401aa161; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_4_io_in_a = io_in_a_4; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_4_io_in_b = 32'h406dd495; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_5_io_in_a = io_in_a_5; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_5_io_in_b = 32'h4060a71d; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_6_io_in_a = io_in_a_6; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_6_io_in_b = 32'h4096fb7e; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_7_io_in_a = io_in_a_7; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_7_io_in_b = 32'h4085b8ba; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_8_io_in_a = io_in_a_8; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_8_io_in_b = 32'h3f25c28e; // @[FPArithmetic.scala 637:33]
  assign FP_adders_0_io_in_a = FP_multipliers_0_io_out_s; // @[FPArithmetic.scala 655:41]
  assign FP_adders_0_io_in_b = FP_multipliers_1_io_out_s; // @[FPArithmetic.scala 656:41]
  assign FP_adders_1_io_in_a = FP_multipliers_2_io_out_s; // @[FPArithmetic.scala 655:41]
  assign FP_adders_1_io_in_b = FP_multipliers_3_io_out_s; // @[FPArithmetic.scala 656:41]
  assign FP_adders_2_io_in_a = FP_multipliers_4_io_out_s; // @[FPArithmetic.scala 655:41]
  assign FP_adders_2_io_in_b = FP_multipliers_5_io_out_s; // @[FPArithmetic.scala 656:41]
  assign FP_adders_3_io_in_a = FP_multipliers_6_io_out_s; // @[FPArithmetic.scala 655:41]
  assign FP_adders_3_io_in_b = FP_multipliers_7_io_out_s; // @[FPArithmetic.scala 656:41]
  assign FP_adders_4_io_in_a = FP_adders_0_io_out_s; // @[FPArithmetic.scala 681:43]
  assign FP_adders_4_io_in_b = FP_adders_1_io_out_s; // @[FPArithmetic.scala 682:43]
  assign FP_adders_5_io_in_a = FP_adders_2_io_out_s; // @[FPArithmetic.scala 681:43]
  assign FP_adders_5_io_in_b = FP_adders_3_io_out_s; // @[FPArithmetic.scala 682:43]
  assign FP_adders_6_io_in_a = FP_adders_4_io_out_s; // @[FPArithmetic.scala 681:43]
  assign FP_adders_6_io_in_b = FP_adders_5_io_out_s; // @[FPArithmetic.scala 682:43]
  assign FP_adders_7_io_in_a = FP_adders_6_io_out_s; // @[FPArithmetic.scala 691:49]
  assign FP_adders_7_io_in_b = FP_multipliers_8_io_out_s; // @[FPArithmetic.scala 650:42]
endmodule
module MatMult1(
  input  [31:0] io_matA_0,
  input  [31:0] io_matA_1,
  input  [31:0] io_matA_2,
  input  [31:0] io_matA_3,
  input  [31:0] io_matA_4,
  input  [31:0] io_matA_5,
  input  [31:0] io_matA_6,
  input  [31:0] io_matA_7,
  input  [31:0] io_matA_8,
  output [31:0] io_f_mac
);
  wire [31:0] f_adder_io_in_a; // @[MatMult.scala 17:25]
  wire [31:0] f_adder_io_in_b; // @[MatMult.scala 17:25]
  wire [31:0] f_adder_io_out_s; // @[MatMult.scala 17:25]
  wire [31:0] mul_io_in_a_0; // @[MatMult.scala 18:21]
  wire [31:0] mul_io_in_a_1; // @[MatMult.scala 18:21]
  wire [31:0] mul_io_in_a_2; // @[MatMult.scala 18:21]
  wire [31:0] mul_io_in_a_3; // @[MatMult.scala 18:21]
  wire [31:0] mul_io_in_a_4; // @[MatMult.scala 18:21]
  wire [31:0] mul_io_in_a_5; // @[MatMult.scala 18:21]
  wire [31:0] mul_io_in_a_6; // @[MatMult.scala 18:21]
  wire [31:0] mul_io_in_a_7; // @[MatMult.scala 18:21]
  wire [31:0] mul_io_in_a_8; // @[MatMult.scala 18:21]
  wire [31:0] mul_io_out_s; // @[MatMult.scala 18:21]
  FP_adder f_adder ( // @[MatMult.scala 17:25]
    .io_in_a(f_adder_io_in_a),
    .io_in_b(f_adder_io_in_b),
    .io_out_s(f_adder_io_out_s)
  );
  FP_multiply_sum mul ( // @[MatMult.scala 18:21]
    .io_in_a_0(mul_io_in_a_0),
    .io_in_a_1(mul_io_in_a_1),
    .io_in_a_2(mul_io_in_a_2),
    .io_in_a_3(mul_io_in_a_3),
    .io_in_a_4(mul_io_in_a_4),
    .io_in_a_5(mul_io_in_a_5),
    .io_in_a_6(mul_io_in_a_6),
    .io_in_a_7(mul_io_in_a_7),
    .io_in_a_8(mul_io_in_a_8),
    .io_out_s(mul_io_out_s)
  );
  assign io_f_mac = f_adder_io_out_s[31] ? 32'h0 : f_adder_io_out_s; // @[MatMult.scala 26:28 27:16 29:16]
  assign f_adder_io_in_a = 32'h1; // @[MatMult.scala 23:21]
  assign f_adder_io_in_b = mul_io_out_s; // @[MatMult.scala 24:21]
  assign mul_io_in_a_0 = io_matA_0; // @[MatMult.scala 20:22]
  assign mul_io_in_a_1 = io_matA_1; // @[MatMult.scala 20:22]
  assign mul_io_in_a_2 = io_matA_2; // @[MatMult.scala 20:22]
  assign mul_io_in_a_3 = io_matA_3; // @[MatMult.scala 20:22]
  assign mul_io_in_a_4 = io_matA_4; // @[MatMult.scala 20:22]
  assign mul_io_in_a_5 = io_matA_5; // @[MatMult.scala 20:22]
  assign mul_io_in_a_6 = io_matA_6; // @[MatMult.scala 20:22]
  assign mul_io_in_a_7 = io_matA_7; // @[MatMult.scala 20:22]
  assign mul_io_in_a_8 = io_matA_8; // @[MatMult.scala 20:22]
endmodule
module Matrix_Controller(
  output [31:0] io_single_out_0,
  output [31:0] io_single_out_1,
  output [31:0] io_single_out_2,
  output [31:0] io_single_out_3,
  output [31:0] io_single_out_4,
  output [31:0] io_single_out_5,
  output [31:0] io_single_out_6,
  output [31:0] io_single_out_7,
  output [31:0] io_single_out_8,
  output [31:0] io_single_out_9,
  output [31:0] io_single_out_10,
  output [31:0] io_single_out_11,
  output [31:0] io_single_out_12,
  output [31:0] io_single_out_13,
  output [31:0] io_single_out_14,
  output [31:0] io_single_out_15,
  output [31:0] io_single_out_16,
  output [31:0] io_single_out_17,
  output [31:0] io_single_out_18,
  output [31:0] io_single_out_19,
  output [31:0] io_single_out_20,
  output [31:0] io_single_out_21,
  output [31:0] io_single_out_22,
  output [31:0] io_single_out_23,
  output [31:0] io_single_out_24,
  output [31:0] io_single_out_25,
  output [31:0] io_single_out_26,
  output [31:0] io_single_out_27,
  output [31:0] io_single_out_28,
  output [31:0] io_single_out_29,
  output [31:0] io_single_out_30,
  output [31:0] io_single_out_31,
  output [31:0] io_single_out_32,
  output [31:0] io_single_out_33,
  output [31:0] io_single_out_34,
  output [31:0] io_single_out_35,
  output [31:0] io_single_out_36,
  output [31:0] io_single_out_37,
  output [31:0] io_single_out_38,
  output [31:0] io_single_out_39,
  output [31:0] io_single_out_40,
  output [31:0] io_single_out_41,
  output [31:0] io_single_out_42,
  output [31:0] io_single_out_43,
  output [31:0] io_single_out_44,
  output [31:0] io_single_out_45,
  output [31:0] io_single_out_46,
  output [31:0] io_single_out_47,
  output [31:0] io_single_out_48,
  output [31:0] io_single_out_49,
  output [31:0] io_single_out_50,
  output [31:0] io_single_out_51,
  output [31:0] io_single_out_52,
  output [31:0] io_single_out_53,
  output [31:0] io_single_out_54,
  output [31:0] io_single_out_55,
  output [31:0] io_single_out_56,
  output [31:0] io_single_out_57,
  output [31:0] io_single_out_58,
  output [31:0] io_single_out_59,
  output [31:0] io_single_out_60,
  output [31:0] io_single_out_61,
  output [31:0] io_single_out_62,
  output [31:0] io_single_out_63
);
  wire [31:0] MatrixMuls_0_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_0_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_0_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_0_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_0_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_0_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_0_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_0_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_0_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_0_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_1_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_1_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_1_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_1_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_1_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_1_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_1_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_1_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_1_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_1_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_2_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_2_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_2_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_2_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_2_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_2_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_2_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_2_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_2_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_2_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_3_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_3_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_3_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_3_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_3_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_3_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_3_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_3_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_3_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_3_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_4_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_4_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_4_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_4_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_4_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_4_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_4_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_4_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_4_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_4_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_5_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_5_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_5_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_5_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_5_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_5_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_5_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_5_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_5_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_5_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_6_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_6_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_6_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_6_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_6_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_6_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_6_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_6_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_6_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_6_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_7_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_7_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_7_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_7_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_7_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_7_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_7_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_7_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_7_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_7_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_8_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_8_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_8_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_8_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_8_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_8_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_8_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_8_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_8_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_8_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_9_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_9_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_9_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_9_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_9_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_9_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_9_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_9_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_9_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_9_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_10_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_10_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_10_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_10_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_10_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_10_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_10_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_10_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_10_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_10_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_11_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_11_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_11_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_11_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_11_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_11_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_11_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_11_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_11_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_11_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_12_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_12_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_12_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_12_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_12_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_12_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_12_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_12_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_12_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_12_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_13_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_13_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_13_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_13_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_13_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_13_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_13_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_13_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_13_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_13_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_14_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_14_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_14_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_14_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_14_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_14_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_14_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_14_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_14_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_14_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_15_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_15_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_15_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_15_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_15_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_15_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_15_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_15_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_15_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_15_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_16_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_16_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_16_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_16_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_16_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_16_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_16_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_16_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_16_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_16_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_17_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_17_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_17_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_17_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_17_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_17_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_17_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_17_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_17_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_17_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_18_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_18_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_18_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_18_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_18_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_18_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_18_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_18_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_18_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_18_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_19_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_19_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_19_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_19_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_19_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_19_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_19_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_19_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_19_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_19_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_20_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_20_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_20_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_20_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_20_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_20_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_20_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_20_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_20_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_20_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_21_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_21_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_21_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_21_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_21_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_21_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_21_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_21_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_21_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_21_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_22_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_22_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_22_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_22_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_22_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_22_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_22_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_22_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_22_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_22_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_23_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_23_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_23_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_23_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_23_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_23_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_23_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_23_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_23_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_23_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_24_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_24_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_24_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_24_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_24_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_24_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_24_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_24_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_24_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_24_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_25_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_25_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_25_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_25_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_25_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_25_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_25_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_25_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_25_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_25_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_26_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_26_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_26_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_26_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_26_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_26_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_26_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_26_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_26_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_26_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_27_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_27_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_27_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_27_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_27_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_27_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_27_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_27_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_27_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_27_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_28_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_28_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_28_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_28_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_28_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_28_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_28_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_28_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_28_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_28_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_29_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_29_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_29_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_29_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_29_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_29_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_29_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_29_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_29_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_29_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_30_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_30_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_30_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_30_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_30_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_30_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_30_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_30_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_30_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_30_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_31_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_31_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_31_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_31_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_31_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_31_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_31_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_31_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_31_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_31_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_32_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_32_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_32_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_32_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_32_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_32_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_32_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_32_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_32_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_32_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_33_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_33_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_33_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_33_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_33_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_33_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_33_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_33_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_33_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_33_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_34_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_34_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_34_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_34_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_34_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_34_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_34_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_34_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_34_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_34_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_35_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_35_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_35_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_35_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_35_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_35_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_35_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_35_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_35_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_35_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_36_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_36_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_36_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_36_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_36_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_36_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_36_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_36_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_36_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_36_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_37_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_37_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_37_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_37_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_37_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_37_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_37_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_37_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_37_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_37_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_38_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_38_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_38_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_38_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_38_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_38_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_38_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_38_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_38_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_38_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_39_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_39_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_39_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_39_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_39_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_39_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_39_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_39_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_39_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_39_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_40_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_40_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_40_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_40_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_40_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_40_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_40_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_40_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_40_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_40_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_41_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_41_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_41_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_41_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_41_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_41_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_41_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_41_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_41_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_41_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_42_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_42_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_42_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_42_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_42_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_42_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_42_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_42_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_42_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_42_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_43_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_43_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_43_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_43_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_43_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_43_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_43_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_43_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_43_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_43_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_44_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_44_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_44_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_44_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_44_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_44_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_44_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_44_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_44_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_44_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_45_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_45_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_45_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_45_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_45_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_45_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_45_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_45_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_45_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_45_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_46_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_46_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_46_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_46_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_46_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_46_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_46_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_46_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_46_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_46_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_47_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_47_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_47_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_47_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_47_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_47_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_47_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_47_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_47_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_47_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_48_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_48_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_48_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_48_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_48_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_48_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_48_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_48_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_48_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_48_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_49_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_49_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_49_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_49_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_49_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_49_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_49_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_49_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_49_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_49_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_50_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_50_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_50_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_50_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_50_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_50_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_50_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_50_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_50_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_50_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_51_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_51_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_51_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_51_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_51_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_51_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_51_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_51_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_51_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_51_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_52_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_52_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_52_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_52_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_52_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_52_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_52_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_52_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_52_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_52_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_53_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_53_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_53_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_53_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_53_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_53_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_53_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_53_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_53_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_53_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_54_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_54_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_54_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_54_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_54_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_54_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_54_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_54_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_54_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_54_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_55_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_55_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_55_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_55_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_55_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_55_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_55_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_55_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_55_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_55_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_56_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_56_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_56_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_56_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_56_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_56_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_56_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_56_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_56_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_56_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_57_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_57_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_57_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_57_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_57_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_57_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_57_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_57_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_57_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_57_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_58_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_58_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_58_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_58_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_58_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_58_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_58_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_58_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_58_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_58_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_59_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_59_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_59_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_59_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_59_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_59_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_59_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_59_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_59_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_59_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_60_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_60_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_60_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_60_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_60_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_60_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_60_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_60_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_60_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_60_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_61_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_61_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_61_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_61_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_61_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_61_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_61_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_61_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_61_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_61_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_62_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_62_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_62_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_62_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_62_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_62_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_62_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_62_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_62_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_62_io_f_mac; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_63_io_matA_0; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_63_io_matA_1; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_63_io_matA_2; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_63_io_matA_3; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_63_io_matA_4; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_63_io_matA_5; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_63_io_matA_6; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_63_io_matA_7; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_63_io_matA_8; // @[Convolution.scala 25:29]
  wire [31:0] MatrixMuls_63_io_f_mac; // @[Convolution.scala 25:29]
  MatMult1 MatrixMuls_0 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_0_io_matA_0),
    .io_matA_1(MatrixMuls_0_io_matA_1),
    .io_matA_2(MatrixMuls_0_io_matA_2),
    .io_matA_3(MatrixMuls_0_io_matA_3),
    .io_matA_4(MatrixMuls_0_io_matA_4),
    .io_matA_5(MatrixMuls_0_io_matA_5),
    .io_matA_6(MatrixMuls_0_io_matA_6),
    .io_matA_7(MatrixMuls_0_io_matA_7),
    .io_matA_8(MatrixMuls_0_io_matA_8),
    .io_f_mac(MatrixMuls_0_io_f_mac)
  );
  MatMult1 MatrixMuls_1 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_1_io_matA_0),
    .io_matA_1(MatrixMuls_1_io_matA_1),
    .io_matA_2(MatrixMuls_1_io_matA_2),
    .io_matA_3(MatrixMuls_1_io_matA_3),
    .io_matA_4(MatrixMuls_1_io_matA_4),
    .io_matA_5(MatrixMuls_1_io_matA_5),
    .io_matA_6(MatrixMuls_1_io_matA_6),
    .io_matA_7(MatrixMuls_1_io_matA_7),
    .io_matA_8(MatrixMuls_1_io_matA_8),
    .io_f_mac(MatrixMuls_1_io_f_mac)
  );
  MatMult1 MatrixMuls_2 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_2_io_matA_0),
    .io_matA_1(MatrixMuls_2_io_matA_1),
    .io_matA_2(MatrixMuls_2_io_matA_2),
    .io_matA_3(MatrixMuls_2_io_matA_3),
    .io_matA_4(MatrixMuls_2_io_matA_4),
    .io_matA_5(MatrixMuls_2_io_matA_5),
    .io_matA_6(MatrixMuls_2_io_matA_6),
    .io_matA_7(MatrixMuls_2_io_matA_7),
    .io_matA_8(MatrixMuls_2_io_matA_8),
    .io_f_mac(MatrixMuls_2_io_f_mac)
  );
  MatMult1 MatrixMuls_3 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_3_io_matA_0),
    .io_matA_1(MatrixMuls_3_io_matA_1),
    .io_matA_2(MatrixMuls_3_io_matA_2),
    .io_matA_3(MatrixMuls_3_io_matA_3),
    .io_matA_4(MatrixMuls_3_io_matA_4),
    .io_matA_5(MatrixMuls_3_io_matA_5),
    .io_matA_6(MatrixMuls_3_io_matA_6),
    .io_matA_7(MatrixMuls_3_io_matA_7),
    .io_matA_8(MatrixMuls_3_io_matA_8),
    .io_f_mac(MatrixMuls_3_io_f_mac)
  );
  MatMult1 MatrixMuls_4 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_4_io_matA_0),
    .io_matA_1(MatrixMuls_4_io_matA_1),
    .io_matA_2(MatrixMuls_4_io_matA_2),
    .io_matA_3(MatrixMuls_4_io_matA_3),
    .io_matA_4(MatrixMuls_4_io_matA_4),
    .io_matA_5(MatrixMuls_4_io_matA_5),
    .io_matA_6(MatrixMuls_4_io_matA_6),
    .io_matA_7(MatrixMuls_4_io_matA_7),
    .io_matA_8(MatrixMuls_4_io_matA_8),
    .io_f_mac(MatrixMuls_4_io_f_mac)
  );
  MatMult1 MatrixMuls_5 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_5_io_matA_0),
    .io_matA_1(MatrixMuls_5_io_matA_1),
    .io_matA_2(MatrixMuls_5_io_matA_2),
    .io_matA_3(MatrixMuls_5_io_matA_3),
    .io_matA_4(MatrixMuls_5_io_matA_4),
    .io_matA_5(MatrixMuls_5_io_matA_5),
    .io_matA_6(MatrixMuls_5_io_matA_6),
    .io_matA_7(MatrixMuls_5_io_matA_7),
    .io_matA_8(MatrixMuls_5_io_matA_8),
    .io_f_mac(MatrixMuls_5_io_f_mac)
  );
  MatMult1 MatrixMuls_6 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_6_io_matA_0),
    .io_matA_1(MatrixMuls_6_io_matA_1),
    .io_matA_2(MatrixMuls_6_io_matA_2),
    .io_matA_3(MatrixMuls_6_io_matA_3),
    .io_matA_4(MatrixMuls_6_io_matA_4),
    .io_matA_5(MatrixMuls_6_io_matA_5),
    .io_matA_6(MatrixMuls_6_io_matA_6),
    .io_matA_7(MatrixMuls_6_io_matA_7),
    .io_matA_8(MatrixMuls_6_io_matA_8),
    .io_f_mac(MatrixMuls_6_io_f_mac)
  );
  MatMult1 MatrixMuls_7 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_7_io_matA_0),
    .io_matA_1(MatrixMuls_7_io_matA_1),
    .io_matA_2(MatrixMuls_7_io_matA_2),
    .io_matA_3(MatrixMuls_7_io_matA_3),
    .io_matA_4(MatrixMuls_7_io_matA_4),
    .io_matA_5(MatrixMuls_7_io_matA_5),
    .io_matA_6(MatrixMuls_7_io_matA_6),
    .io_matA_7(MatrixMuls_7_io_matA_7),
    .io_matA_8(MatrixMuls_7_io_matA_8),
    .io_f_mac(MatrixMuls_7_io_f_mac)
  );
  MatMult1 MatrixMuls_8 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_8_io_matA_0),
    .io_matA_1(MatrixMuls_8_io_matA_1),
    .io_matA_2(MatrixMuls_8_io_matA_2),
    .io_matA_3(MatrixMuls_8_io_matA_3),
    .io_matA_4(MatrixMuls_8_io_matA_4),
    .io_matA_5(MatrixMuls_8_io_matA_5),
    .io_matA_6(MatrixMuls_8_io_matA_6),
    .io_matA_7(MatrixMuls_8_io_matA_7),
    .io_matA_8(MatrixMuls_8_io_matA_8),
    .io_f_mac(MatrixMuls_8_io_f_mac)
  );
  MatMult1 MatrixMuls_9 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_9_io_matA_0),
    .io_matA_1(MatrixMuls_9_io_matA_1),
    .io_matA_2(MatrixMuls_9_io_matA_2),
    .io_matA_3(MatrixMuls_9_io_matA_3),
    .io_matA_4(MatrixMuls_9_io_matA_4),
    .io_matA_5(MatrixMuls_9_io_matA_5),
    .io_matA_6(MatrixMuls_9_io_matA_6),
    .io_matA_7(MatrixMuls_9_io_matA_7),
    .io_matA_8(MatrixMuls_9_io_matA_8),
    .io_f_mac(MatrixMuls_9_io_f_mac)
  );
  MatMult1 MatrixMuls_10 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_10_io_matA_0),
    .io_matA_1(MatrixMuls_10_io_matA_1),
    .io_matA_2(MatrixMuls_10_io_matA_2),
    .io_matA_3(MatrixMuls_10_io_matA_3),
    .io_matA_4(MatrixMuls_10_io_matA_4),
    .io_matA_5(MatrixMuls_10_io_matA_5),
    .io_matA_6(MatrixMuls_10_io_matA_6),
    .io_matA_7(MatrixMuls_10_io_matA_7),
    .io_matA_8(MatrixMuls_10_io_matA_8),
    .io_f_mac(MatrixMuls_10_io_f_mac)
  );
  MatMult1 MatrixMuls_11 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_11_io_matA_0),
    .io_matA_1(MatrixMuls_11_io_matA_1),
    .io_matA_2(MatrixMuls_11_io_matA_2),
    .io_matA_3(MatrixMuls_11_io_matA_3),
    .io_matA_4(MatrixMuls_11_io_matA_4),
    .io_matA_5(MatrixMuls_11_io_matA_5),
    .io_matA_6(MatrixMuls_11_io_matA_6),
    .io_matA_7(MatrixMuls_11_io_matA_7),
    .io_matA_8(MatrixMuls_11_io_matA_8),
    .io_f_mac(MatrixMuls_11_io_f_mac)
  );
  MatMult1 MatrixMuls_12 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_12_io_matA_0),
    .io_matA_1(MatrixMuls_12_io_matA_1),
    .io_matA_2(MatrixMuls_12_io_matA_2),
    .io_matA_3(MatrixMuls_12_io_matA_3),
    .io_matA_4(MatrixMuls_12_io_matA_4),
    .io_matA_5(MatrixMuls_12_io_matA_5),
    .io_matA_6(MatrixMuls_12_io_matA_6),
    .io_matA_7(MatrixMuls_12_io_matA_7),
    .io_matA_8(MatrixMuls_12_io_matA_8),
    .io_f_mac(MatrixMuls_12_io_f_mac)
  );
  MatMult1 MatrixMuls_13 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_13_io_matA_0),
    .io_matA_1(MatrixMuls_13_io_matA_1),
    .io_matA_2(MatrixMuls_13_io_matA_2),
    .io_matA_3(MatrixMuls_13_io_matA_3),
    .io_matA_4(MatrixMuls_13_io_matA_4),
    .io_matA_5(MatrixMuls_13_io_matA_5),
    .io_matA_6(MatrixMuls_13_io_matA_6),
    .io_matA_7(MatrixMuls_13_io_matA_7),
    .io_matA_8(MatrixMuls_13_io_matA_8),
    .io_f_mac(MatrixMuls_13_io_f_mac)
  );
  MatMult1 MatrixMuls_14 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_14_io_matA_0),
    .io_matA_1(MatrixMuls_14_io_matA_1),
    .io_matA_2(MatrixMuls_14_io_matA_2),
    .io_matA_3(MatrixMuls_14_io_matA_3),
    .io_matA_4(MatrixMuls_14_io_matA_4),
    .io_matA_5(MatrixMuls_14_io_matA_5),
    .io_matA_6(MatrixMuls_14_io_matA_6),
    .io_matA_7(MatrixMuls_14_io_matA_7),
    .io_matA_8(MatrixMuls_14_io_matA_8),
    .io_f_mac(MatrixMuls_14_io_f_mac)
  );
  MatMult1 MatrixMuls_15 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_15_io_matA_0),
    .io_matA_1(MatrixMuls_15_io_matA_1),
    .io_matA_2(MatrixMuls_15_io_matA_2),
    .io_matA_3(MatrixMuls_15_io_matA_3),
    .io_matA_4(MatrixMuls_15_io_matA_4),
    .io_matA_5(MatrixMuls_15_io_matA_5),
    .io_matA_6(MatrixMuls_15_io_matA_6),
    .io_matA_7(MatrixMuls_15_io_matA_7),
    .io_matA_8(MatrixMuls_15_io_matA_8),
    .io_f_mac(MatrixMuls_15_io_f_mac)
  );
  MatMult1 MatrixMuls_16 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_16_io_matA_0),
    .io_matA_1(MatrixMuls_16_io_matA_1),
    .io_matA_2(MatrixMuls_16_io_matA_2),
    .io_matA_3(MatrixMuls_16_io_matA_3),
    .io_matA_4(MatrixMuls_16_io_matA_4),
    .io_matA_5(MatrixMuls_16_io_matA_5),
    .io_matA_6(MatrixMuls_16_io_matA_6),
    .io_matA_7(MatrixMuls_16_io_matA_7),
    .io_matA_8(MatrixMuls_16_io_matA_8),
    .io_f_mac(MatrixMuls_16_io_f_mac)
  );
  MatMult1 MatrixMuls_17 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_17_io_matA_0),
    .io_matA_1(MatrixMuls_17_io_matA_1),
    .io_matA_2(MatrixMuls_17_io_matA_2),
    .io_matA_3(MatrixMuls_17_io_matA_3),
    .io_matA_4(MatrixMuls_17_io_matA_4),
    .io_matA_5(MatrixMuls_17_io_matA_5),
    .io_matA_6(MatrixMuls_17_io_matA_6),
    .io_matA_7(MatrixMuls_17_io_matA_7),
    .io_matA_8(MatrixMuls_17_io_matA_8),
    .io_f_mac(MatrixMuls_17_io_f_mac)
  );
  MatMult1 MatrixMuls_18 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_18_io_matA_0),
    .io_matA_1(MatrixMuls_18_io_matA_1),
    .io_matA_2(MatrixMuls_18_io_matA_2),
    .io_matA_3(MatrixMuls_18_io_matA_3),
    .io_matA_4(MatrixMuls_18_io_matA_4),
    .io_matA_5(MatrixMuls_18_io_matA_5),
    .io_matA_6(MatrixMuls_18_io_matA_6),
    .io_matA_7(MatrixMuls_18_io_matA_7),
    .io_matA_8(MatrixMuls_18_io_matA_8),
    .io_f_mac(MatrixMuls_18_io_f_mac)
  );
  MatMult1 MatrixMuls_19 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_19_io_matA_0),
    .io_matA_1(MatrixMuls_19_io_matA_1),
    .io_matA_2(MatrixMuls_19_io_matA_2),
    .io_matA_3(MatrixMuls_19_io_matA_3),
    .io_matA_4(MatrixMuls_19_io_matA_4),
    .io_matA_5(MatrixMuls_19_io_matA_5),
    .io_matA_6(MatrixMuls_19_io_matA_6),
    .io_matA_7(MatrixMuls_19_io_matA_7),
    .io_matA_8(MatrixMuls_19_io_matA_8),
    .io_f_mac(MatrixMuls_19_io_f_mac)
  );
  MatMult1 MatrixMuls_20 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_20_io_matA_0),
    .io_matA_1(MatrixMuls_20_io_matA_1),
    .io_matA_2(MatrixMuls_20_io_matA_2),
    .io_matA_3(MatrixMuls_20_io_matA_3),
    .io_matA_4(MatrixMuls_20_io_matA_4),
    .io_matA_5(MatrixMuls_20_io_matA_5),
    .io_matA_6(MatrixMuls_20_io_matA_6),
    .io_matA_7(MatrixMuls_20_io_matA_7),
    .io_matA_8(MatrixMuls_20_io_matA_8),
    .io_f_mac(MatrixMuls_20_io_f_mac)
  );
  MatMult1 MatrixMuls_21 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_21_io_matA_0),
    .io_matA_1(MatrixMuls_21_io_matA_1),
    .io_matA_2(MatrixMuls_21_io_matA_2),
    .io_matA_3(MatrixMuls_21_io_matA_3),
    .io_matA_4(MatrixMuls_21_io_matA_4),
    .io_matA_5(MatrixMuls_21_io_matA_5),
    .io_matA_6(MatrixMuls_21_io_matA_6),
    .io_matA_7(MatrixMuls_21_io_matA_7),
    .io_matA_8(MatrixMuls_21_io_matA_8),
    .io_f_mac(MatrixMuls_21_io_f_mac)
  );
  MatMult1 MatrixMuls_22 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_22_io_matA_0),
    .io_matA_1(MatrixMuls_22_io_matA_1),
    .io_matA_2(MatrixMuls_22_io_matA_2),
    .io_matA_3(MatrixMuls_22_io_matA_3),
    .io_matA_4(MatrixMuls_22_io_matA_4),
    .io_matA_5(MatrixMuls_22_io_matA_5),
    .io_matA_6(MatrixMuls_22_io_matA_6),
    .io_matA_7(MatrixMuls_22_io_matA_7),
    .io_matA_8(MatrixMuls_22_io_matA_8),
    .io_f_mac(MatrixMuls_22_io_f_mac)
  );
  MatMult1 MatrixMuls_23 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_23_io_matA_0),
    .io_matA_1(MatrixMuls_23_io_matA_1),
    .io_matA_2(MatrixMuls_23_io_matA_2),
    .io_matA_3(MatrixMuls_23_io_matA_3),
    .io_matA_4(MatrixMuls_23_io_matA_4),
    .io_matA_5(MatrixMuls_23_io_matA_5),
    .io_matA_6(MatrixMuls_23_io_matA_6),
    .io_matA_7(MatrixMuls_23_io_matA_7),
    .io_matA_8(MatrixMuls_23_io_matA_8),
    .io_f_mac(MatrixMuls_23_io_f_mac)
  );
  MatMult1 MatrixMuls_24 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_24_io_matA_0),
    .io_matA_1(MatrixMuls_24_io_matA_1),
    .io_matA_2(MatrixMuls_24_io_matA_2),
    .io_matA_3(MatrixMuls_24_io_matA_3),
    .io_matA_4(MatrixMuls_24_io_matA_4),
    .io_matA_5(MatrixMuls_24_io_matA_5),
    .io_matA_6(MatrixMuls_24_io_matA_6),
    .io_matA_7(MatrixMuls_24_io_matA_7),
    .io_matA_8(MatrixMuls_24_io_matA_8),
    .io_f_mac(MatrixMuls_24_io_f_mac)
  );
  MatMult1 MatrixMuls_25 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_25_io_matA_0),
    .io_matA_1(MatrixMuls_25_io_matA_1),
    .io_matA_2(MatrixMuls_25_io_matA_2),
    .io_matA_3(MatrixMuls_25_io_matA_3),
    .io_matA_4(MatrixMuls_25_io_matA_4),
    .io_matA_5(MatrixMuls_25_io_matA_5),
    .io_matA_6(MatrixMuls_25_io_matA_6),
    .io_matA_7(MatrixMuls_25_io_matA_7),
    .io_matA_8(MatrixMuls_25_io_matA_8),
    .io_f_mac(MatrixMuls_25_io_f_mac)
  );
  MatMult1 MatrixMuls_26 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_26_io_matA_0),
    .io_matA_1(MatrixMuls_26_io_matA_1),
    .io_matA_2(MatrixMuls_26_io_matA_2),
    .io_matA_3(MatrixMuls_26_io_matA_3),
    .io_matA_4(MatrixMuls_26_io_matA_4),
    .io_matA_5(MatrixMuls_26_io_matA_5),
    .io_matA_6(MatrixMuls_26_io_matA_6),
    .io_matA_7(MatrixMuls_26_io_matA_7),
    .io_matA_8(MatrixMuls_26_io_matA_8),
    .io_f_mac(MatrixMuls_26_io_f_mac)
  );
  MatMult1 MatrixMuls_27 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_27_io_matA_0),
    .io_matA_1(MatrixMuls_27_io_matA_1),
    .io_matA_2(MatrixMuls_27_io_matA_2),
    .io_matA_3(MatrixMuls_27_io_matA_3),
    .io_matA_4(MatrixMuls_27_io_matA_4),
    .io_matA_5(MatrixMuls_27_io_matA_5),
    .io_matA_6(MatrixMuls_27_io_matA_6),
    .io_matA_7(MatrixMuls_27_io_matA_7),
    .io_matA_8(MatrixMuls_27_io_matA_8),
    .io_f_mac(MatrixMuls_27_io_f_mac)
  );
  MatMult1 MatrixMuls_28 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_28_io_matA_0),
    .io_matA_1(MatrixMuls_28_io_matA_1),
    .io_matA_2(MatrixMuls_28_io_matA_2),
    .io_matA_3(MatrixMuls_28_io_matA_3),
    .io_matA_4(MatrixMuls_28_io_matA_4),
    .io_matA_5(MatrixMuls_28_io_matA_5),
    .io_matA_6(MatrixMuls_28_io_matA_6),
    .io_matA_7(MatrixMuls_28_io_matA_7),
    .io_matA_8(MatrixMuls_28_io_matA_8),
    .io_f_mac(MatrixMuls_28_io_f_mac)
  );
  MatMult1 MatrixMuls_29 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_29_io_matA_0),
    .io_matA_1(MatrixMuls_29_io_matA_1),
    .io_matA_2(MatrixMuls_29_io_matA_2),
    .io_matA_3(MatrixMuls_29_io_matA_3),
    .io_matA_4(MatrixMuls_29_io_matA_4),
    .io_matA_5(MatrixMuls_29_io_matA_5),
    .io_matA_6(MatrixMuls_29_io_matA_6),
    .io_matA_7(MatrixMuls_29_io_matA_7),
    .io_matA_8(MatrixMuls_29_io_matA_8),
    .io_f_mac(MatrixMuls_29_io_f_mac)
  );
  MatMult1 MatrixMuls_30 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_30_io_matA_0),
    .io_matA_1(MatrixMuls_30_io_matA_1),
    .io_matA_2(MatrixMuls_30_io_matA_2),
    .io_matA_3(MatrixMuls_30_io_matA_3),
    .io_matA_4(MatrixMuls_30_io_matA_4),
    .io_matA_5(MatrixMuls_30_io_matA_5),
    .io_matA_6(MatrixMuls_30_io_matA_6),
    .io_matA_7(MatrixMuls_30_io_matA_7),
    .io_matA_8(MatrixMuls_30_io_matA_8),
    .io_f_mac(MatrixMuls_30_io_f_mac)
  );
  MatMult1 MatrixMuls_31 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_31_io_matA_0),
    .io_matA_1(MatrixMuls_31_io_matA_1),
    .io_matA_2(MatrixMuls_31_io_matA_2),
    .io_matA_3(MatrixMuls_31_io_matA_3),
    .io_matA_4(MatrixMuls_31_io_matA_4),
    .io_matA_5(MatrixMuls_31_io_matA_5),
    .io_matA_6(MatrixMuls_31_io_matA_6),
    .io_matA_7(MatrixMuls_31_io_matA_7),
    .io_matA_8(MatrixMuls_31_io_matA_8),
    .io_f_mac(MatrixMuls_31_io_f_mac)
  );
  MatMult1 MatrixMuls_32 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_32_io_matA_0),
    .io_matA_1(MatrixMuls_32_io_matA_1),
    .io_matA_2(MatrixMuls_32_io_matA_2),
    .io_matA_3(MatrixMuls_32_io_matA_3),
    .io_matA_4(MatrixMuls_32_io_matA_4),
    .io_matA_5(MatrixMuls_32_io_matA_5),
    .io_matA_6(MatrixMuls_32_io_matA_6),
    .io_matA_7(MatrixMuls_32_io_matA_7),
    .io_matA_8(MatrixMuls_32_io_matA_8),
    .io_f_mac(MatrixMuls_32_io_f_mac)
  );
  MatMult1 MatrixMuls_33 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_33_io_matA_0),
    .io_matA_1(MatrixMuls_33_io_matA_1),
    .io_matA_2(MatrixMuls_33_io_matA_2),
    .io_matA_3(MatrixMuls_33_io_matA_3),
    .io_matA_4(MatrixMuls_33_io_matA_4),
    .io_matA_5(MatrixMuls_33_io_matA_5),
    .io_matA_6(MatrixMuls_33_io_matA_6),
    .io_matA_7(MatrixMuls_33_io_matA_7),
    .io_matA_8(MatrixMuls_33_io_matA_8),
    .io_f_mac(MatrixMuls_33_io_f_mac)
  );
  MatMult1 MatrixMuls_34 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_34_io_matA_0),
    .io_matA_1(MatrixMuls_34_io_matA_1),
    .io_matA_2(MatrixMuls_34_io_matA_2),
    .io_matA_3(MatrixMuls_34_io_matA_3),
    .io_matA_4(MatrixMuls_34_io_matA_4),
    .io_matA_5(MatrixMuls_34_io_matA_5),
    .io_matA_6(MatrixMuls_34_io_matA_6),
    .io_matA_7(MatrixMuls_34_io_matA_7),
    .io_matA_8(MatrixMuls_34_io_matA_8),
    .io_f_mac(MatrixMuls_34_io_f_mac)
  );
  MatMult1 MatrixMuls_35 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_35_io_matA_0),
    .io_matA_1(MatrixMuls_35_io_matA_1),
    .io_matA_2(MatrixMuls_35_io_matA_2),
    .io_matA_3(MatrixMuls_35_io_matA_3),
    .io_matA_4(MatrixMuls_35_io_matA_4),
    .io_matA_5(MatrixMuls_35_io_matA_5),
    .io_matA_6(MatrixMuls_35_io_matA_6),
    .io_matA_7(MatrixMuls_35_io_matA_7),
    .io_matA_8(MatrixMuls_35_io_matA_8),
    .io_f_mac(MatrixMuls_35_io_f_mac)
  );
  MatMult1 MatrixMuls_36 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_36_io_matA_0),
    .io_matA_1(MatrixMuls_36_io_matA_1),
    .io_matA_2(MatrixMuls_36_io_matA_2),
    .io_matA_3(MatrixMuls_36_io_matA_3),
    .io_matA_4(MatrixMuls_36_io_matA_4),
    .io_matA_5(MatrixMuls_36_io_matA_5),
    .io_matA_6(MatrixMuls_36_io_matA_6),
    .io_matA_7(MatrixMuls_36_io_matA_7),
    .io_matA_8(MatrixMuls_36_io_matA_8),
    .io_f_mac(MatrixMuls_36_io_f_mac)
  );
  MatMult1 MatrixMuls_37 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_37_io_matA_0),
    .io_matA_1(MatrixMuls_37_io_matA_1),
    .io_matA_2(MatrixMuls_37_io_matA_2),
    .io_matA_3(MatrixMuls_37_io_matA_3),
    .io_matA_4(MatrixMuls_37_io_matA_4),
    .io_matA_5(MatrixMuls_37_io_matA_5),
    .io_matA_6(MatrixMuls_37_io_matA_6),
    .io_matA_7(MatrixMuls_37_io_matA_7),
    .io_matA_8(MatrixMuls_37_io_matA_8),
    .io_f_mac(MatrixMuls_37_io_f_mac)
  );
  MatMult1 MatrixMuls_38 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_38_io_matA_0),
    .io_matA_1(MatrixMuls_38_io_matA_1),
    .io_matA_2(MatrixMuls_38_io_matA_2),
    .io_matA_3(MatrixMuls_38_io_matA_3),
    .io_matA_4(MatrixMuls_38_io_matA_4),
    .io_matA_5(MatrixMuls_38_io_matA_5),
    .io_matA_6(MatrixMuls_38_io_matA_6),
    .io_matA_7(MatrixMuls_38_io_matA_7),
    .io_matA_8(MatrixMuls_38_io_matA_8),
    .io_f_mac(MatrixMuls_38_io_f_mac)
  );
  MatMult1 MatrixMuls_39 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_39_io_matA_0),
    .io_matA_1(MatrixMuls_39_io_matA_1),
    .io_matA_2(MatrixMuls_39_io_matA_2),
    .io_matA_3(MatrixMuls_39_io_matA_3),
    .io_matA_4(MatrixMuls_39_io_matA_4),
    .io_matA_5(MatrixMuls_39_io_matA_5),
    .io_matA_6(MatrixMuls_39_io_matA_6),
    .io_matA_7(MatrixMuls_39_io_matA_7),
    .io_matA_8(MatrixMuls_39_io_matA_8),
    .io_f_mac(MatrixMuls_39_io_f_mac)
  );
  MatMult1 MatrixMuls_40 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_40_io_matA_0),
    .io_matA_1(MatrixMuls_40_io_matA_1),
    .io_matA_2(MatrixMuls_40_io_matA_2),
    .io_matA_3(MatrixMuls_40_io_matA_3),
    .io_matA_4(MatrixMuls_40_io_matA_4),
    .io_matA_5(MatrixMuls_40_io_matA_5),
    .io_matA_6(MatrixMuls_40_io_matA_6),
    .io_matA_7(MatrixMuls_40_io_matA_7),
    .io_matA_8(MatrixMuls_40_io_matA_8),
    .io_f_mac(MatrixMuls_40_io_f_mac)
  );
  MatMult1 MatrixMuls_41 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_41_io_matA_0),
    .io_matA_1(MatrixMuls_41_io_matA_1),
    .io_matA_2(MatrixMuls_41_io_matA_2),
    .io_matA_3(MatrixMuls_41_io_matA_3),
    .io_matA_4(MatrixMuls_41_io_matA_4),
    .io_matA_5(MatrixMuls_41_io_matA_5),
    .io_matA_6(MatrixMuls_41_io_matA_6),
    .io_matA_7(MatrixMuls_41_io_matA_7),
    .io_matA_8(MatrixMuls_41_io_matA_8),
    .io_f_mac(MatrixMuls_41_io_f_mac)
  );
  MatMult1 MatrixMuls_42 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_42_io_matA_0),
    .io_matA_1(MatrixMuls_42_io_matA_1),
    .io_matA_2(MatrixMuls_42_io_matA_2),
    .io_matA_3(MatrixMuls_42_io_matA_3),
    .io_matA_4(MatrixMuls_42_io_matA_4),
    .io_matA_5(MatrixMuls_42_io_matA_5),
    .io_matA_6(MatrixMuls_42_io_matA_6),
    .io_matA_7(MatrixMuls_42_io_matA_7),
    .io_matA_8(MatrixMuls_42_io_matA_8),
    .io_f_mac(MatrixMuls_42_io_f_mac)
  );
  MatMult1 MatrixMuls_43 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_43_io_matA_0),
    .io_matA_1(MatrixMuls_43_io_matA_1),
    .io_matA_2(MatrixMuls_43_io_matA_2),
    .io_matA_3(MatrixMuls_43_io_matA_3),
    .io_matA_4(MatrixMuls_43_io_matA_4),
    .io_matA_5(MatrixMuls_43_io_matA_5),
    .io_matA_6(MatrixMuls_43_io_matA_6),
    .io_matA_7(MatrixMuls_43_io_matA_7),
    .io_matA_8(MatrixMuls_43_io_matA_8),
    .io_f_mac(MatrixMuls_43_io_f_mac)
  );
  MatMult1 MatrixMuls_44 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_44_io_matA_0),
    .io_matA_1(MatrixMuls_44_io_matA_1),
    .io_matA_2(MatrixMuls_44_io_matA_2),
    .io_matA_3(MatrixMuls_44_io_matA_3),
    .io_matA_4(MatrixMuls_44_io_matA_4),
    .io_matA_5(MatrixMuls_44_io_matA_5),
    .io_matA_6(MatrixMuls_44_io_matA_6),
    .io_matA_7(MatrixMuls_44_io_matA_7),
    .io_matA_8(MatrixMuls_44_io_matA_8),
    .io_f_mac(MatrixMuls_44_io_f_mac)
  );
  MatMult1 MatrixMuls_45 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_45_io_matA_0),
    .io_matA_1(MatrixMuls_45_io_matA_1),
    .io_matA_2(MatrixMuls_45_io_matA_2),
    .io_matA_3(MatrixMuls_45_io_matA_3),
    .io_matA_4(MatrixMuls_45_io_matA_4),
    .io_matA_5(MatrixMuls_45_io_matA_5),
    .io_matA_6(MatrixMuls_45_io_matA_6),
    .io_matA_7(MatrixMuls_45_io_matA_7),
    .io_matA_8(MatrixMuls_45_io_matA_8),
    .io_f_mac(MatrixMuls_45_io_f_mac)
  );
  MatMult1 MatrixMuls_46 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_46_io_matA_0),
    .io_matA_1(MatrixMuls_46_io_matA_1),
    .io_matA_2(MatrixMuls_46_io_matA_2),
    .io_matA_3(MatrixMuls_46_io_matA_3),
    .io_matA_4(MatrixMuls_46_io_matA_4),
    .io_matA_5(MatrixMuls_46_io_matA_5),
    .io_matA_6(MatrixMuls_46_io_matA_6),
    .io_matA_7(MatrixMuls_46_io_matA_7),
    .io_matA_8(MatrixMuls_46_io_matA_8),
    .io_f_mac(MatrixMuls_46_io_f_mac)
  );
  MatMult1 MatrixMuls_47 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_47_io_matA_0),
    .io_matA_1(MatrixMuls_47_io_matA_1),
    .io_matA_2(MatrixMuls_47_io_matA_2),
    .io_matA_3(MatrixMuls_47_io_matA_3),
    .io_matA_4(MatrixMuls_47_io_matA_4),
    .io_matA_5(MatrixMuls_47_io_matA_5),
    .io_matA_6(MatrixMuls_47_io_matA_6),
    .io_matA_7(MatrixMuls_47_io_matA_7),
    .io_matA_8(MatrixMuls_47_io_matA_8),
    .io_f_mac(MatrixMuls_47_io_f_mac)
  );
  MatMult1 MatrixMuls_48 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_48_io_matA_0),
    .io_matA_1(MatrixMuls_48_io_matA_1),
    .io_matA_2(MatrixMuls_48_io_matA_2),
    .io_matA_3(MatrixMuls_48_io_matA_3),
    .io_matA_4(MatrixMuls_48_io_matA_4),
    .io_matA_5(MatrixMuls_48_io_matA_5),
    .io_matA_6(MatrixMuls_48_io_matA_6),
    .io_matA_7(MatrixMuls_48_io_matA_7),
    .io_matA_8(MatrixMuls_48_io_matA_8),
    .io_f_mac(MatrixMuls_48_io_f_mac)
  );
  MatMult1 MatrixMuls_49 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_49_io_matA_0),
    .io_matA_1(MatrixMuls_49_io_matA_1),
    .io_matA_2(MatrixMuls_49_io_matA_2),
    .io_matA_3(MatrixMuls_49_io_matA_3),
    .io_matA_4(MatrixMuls_49_io_matA_4),
    .io_matA_5(MatrixMuls_49_io_matA_5),
    .io_matA_6(MatrixMuls_49_io_matA_6),
    .io_matA_7(MatrixMuls_49_io_matA_7),
    .io_matA_8(MatrixMuls_49_io_matA_8),
    .io_f_mac(MatrixMuls_49_io_f_mac)
  );
  MatMult1 MatrixMuls_50 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_50_io_matA_0),
    .io_matA_1(MatrixMuls_50_io_matA_1),
    .io_matA_2(MatrixMuls_50_io_matA_2),
    .io_matA_3(MatrixMuls_50_io_matA_3),
    .io_matA_4(MatrixMuls_50_io_matA_4),
    .io_matA_5(MatrixMuls_50_io_matA_5),
    .io_matA_6(MatrixMuls_50_io_matA_6),
    .io_matA_7(MatrixMuls_50_io_matA_7),
    .io_matA_8(MatrixMuls_50_io_matA_8),
    .io_f_mac(MatrixMuls_50_io_f_mac)
  );
  MatMult1 MatrixMuls_51 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_51_io_matA_0),
    .io_matA_1(MatrixMuls_51_io_matA_1),
    .io_matA_2(MatrixMuls_51_io_matA_2),
    .io_matA_3(MatrixMuls_51_io_matA_3),
    .io_matA_4(MatrixMuls_51_io_matA_4),
    .io_matA_5(MatrixMuls_51_io_matA_5),
    .io_matA_6(MatrixMuls_51_io_matA_6),
    .io_matA_7(MatrixMuls_51_io_matA_7),
    .io_matA_8(MatrixMuls_51_io_matA_8),
    .io_f_mac(MatrixMuls_51_io_f_mac)
  );
  MatMult1 MatrixMuls_52 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_52_io_matA_0),
    .io_matA_1(MatrixMuls_52_io_matA_1),
    .io_matA_2(MatrixMuls_52_io_matA_2),
    .io_matA_3(MatrixMuls_52_io_matA_3),
    .io_matA_4(MatrixMuls_52_io_matA_4),
    .io_matA_5(MatrixMuls_52_io_matA_5),
    .io_matA_6(MatrixMuls_52_io_matA_6),
    .io_matA_7(MatrixMuls_52_io_matA_7),
    .io_matA_8(MatrixMuls_52_io_matA_8),
    .io_f_mac(MatrixMuls_52_io_f_mac)
  );
  MatMult1 MatrixMuls_53 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_53_io_matA_0),
    .io_matA_1(MatrixMuls_53_io_matA_1),
    .io_matA_2(MatrixMuls_53_io_matA_2),
    .io_matA_3(MatrixMuls_53_io_matA_3),
    .io_matA_4(MatrixMuls_53_io_matA_4),
    .io_matA_5(MatrixMuls_53_io_matA_5),
    .io_matA_6(MatrixMuls_53_io_matA_6),
    .io_matA_7(MatrixMuls_53_io_matA_7),
    .io_matA_8(MatrixMuls_53_io_matA_8),
    .io_f_mac(MatrixMuls_53_io_f_mac)
  );
  MatMult1 MatrixMuls_54 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_54_io_matA_0),
    .io_matA_1(MatrixMuls_54_io_matA_1),
    .io_matA_2(MatrixMuls_54_io_matA_2),
    .io_matA_3(MatrixMuls_54_io_matA_3),
    .io_matA_4(MatrixMuls_54_io_matA_4),
    .io_matA_5(MatrixMuls_54_io_matA_5),
    .io_matA_6(MatrixMuls_54_io_matA_6),
    .io_matA_7(MatrixMuls_54_io_matA_7),
    .io_matA_8(MatrixMuls_54_io_matA_8),
    .io_f_mac(MatrixMuls_54_io_f_mac)
  );
  MatMult1 MatrixMuls_55 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_55_io_matA_0),
    .io_matA_1(MatrixMuls_55_io_matA_1),
    .io_matA_2(MatrixMuls_55_io_matA_2),
    .io_matA_3(MatrixMuls_55_io_matA_3),
    .io_matA_4(MatrixMuls_55_io_matA_4),
    .io_matA_5(MatrixMuls_55_io_matA_5),
    .io_matA_6(MatrixMuls_55_io_matA_6),
    .io_matA_7(MatrixMuls_55_io_matA_7),
    .io_matA_8(MatrixMuls_55_io_matA_8),
    .io_f_mac(MatrixMuls_55_io_f_mac)
  );
  MatMult1 MatrixMuls_56 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_56_io_matA_0),
    .io_matA_1(MatrixMuls_56_io_matA_1),
    .io_matA_2(MatrixMuls_56_io_matA_2),
    .io_matA_3(MatrixMuls_56_io_matA_3),
    .io_matA_4(MatrixMuls_56_io_matA_4),
    .io_matA_5(MatrixMuls_56_io_matA_5),
    .io_matA_6(MatrixMuls_56_io_matA_6),
    .io_matA_7(MatrixMuls_56_io_matA_7),
    .io_matA_8(MatrixMuls_56_io_matA_8),
    .io_f_mac(MatrixMuls_56_io_f_mac)
  );
  MatMult1 MatrixMuls_57 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_57_io_matA_0),
    .io_matA_1(MatrixMuls_57_io_matA_1),
    .io_matA_2(MatrixMuls_57_io_matA_2),
    .io_matA_3(MatrixMuls_57_io_matA_3),
    .io_matA_4(MatrixMuls_57_io_matA_4),
    .io_matA_5(MatrixMuls_57_io_matA_5),
    .io_matA_6(MatrixMuls_57_io_matA_6),
    .io_matA_7(MatrixMuls_57_io_matA_7),
    .io_matA_8(MatrixMuls_57_io_matA_8),
    .io_f_mac(MatrixMuls_57_io_f_mac)
  );
  MatMult1 MatrixMuls_58 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_58_io_matA_0),
    .io_matA_1(MatrixMuls_58_io_matA_1),
    .io_matA_2(MatrixMuls_58_io_matA_2),
    .io_matA_3(MatrixMuls_58_io_matA_3),
    .io_matA_4(MatrixMuls_58_io_matA_4),
    .io_matA_5(MatrixMuls_58_io_matA_5),
    .io_matA_6(MatrixMuls_58_io_matA_6),
    .io_matA_7(MatrixMuls_58_io_matA_7),
    .io_matA_8(MatrixMuls_58_io_matA_8),
    .io_f_mac(MatrixMuls_58_io_f_mac)
  );
  MatMult1 MatrixMuls_59 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_59_io_matA_0),
    .io_matA_1(MatrixMuls_59_io_matA_1),
    .io_matA_2(MatrixMuls_59_io_matA_2),
    .io_matA_3(MatrixMuls_59_io_matA_3),
    .io_matA_4(MatrixMuls_59_io_matA_4),
    .io_matA_5(MatrixMuls_59_io_matA_5),
    .io_matA_6(MatrixMuls_59_io_matA_6),
    .io_matA_7(MatrixMuls_59_io_matA_7),
    .io_matA_8(MatrixMuls_59_io_matA_8),
    .io_f_mac(MatrixMuls_59_io_f_mac)
  );
  MatMult1 MatrixMuls_60 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_60_io_matA_0),
    .io_matA_1(MatrixMuls_60_io_matA_1),
    .io_matA_2(MatrixMuls_60_io_matA_2),
    .io_matA_3(MatrixMuls_60_io_matA_3),
    .io_matA_4(MatrixMuls_60_io_matA_4),
    .io_matA_5(MatrixMuls_60_io_matA_5),
    .io_matA_6(MatrixMuls_60_io_matA_6),
    .io_matA_7(MatrixMuls_60_io_matA_7),
    .io_matA_8(MatrixMuls_60_io_matA_8),
    .io_f_mac(MatrixMuls_60_io_f_mac)
  );
  MatMult1 MatrixMuls_61 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_61_io_matA_0),
    .io_matA_1(MatrixMuls_61_io_matA_1),
    .io_matA_2(MatrixMuls_61_io_matA_2),
    .io_matA_3(MatrixMuls_61_io_matA_3),
    .io_matA_4(MatrixMuls_61_io_matA_4),
    .io_matA_5(MatrixMuls_61_io_matA_5),
    .io_matA_6(MatrixMuls_61_io_matA_6),
    .io_matA_7(MatrixMuls_61_io_matA_7),
    .io_matA_8(MatrixMuls_61_io_matA_8),
    .io_f_mac(MatrixMuls_61_io_f_mac)
  );
  MatMult1 MatrixMuls_62 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_62_io_matA_0),
    .io_matA_1(MatrixMuls_62_io_matA_1),
    .io_matA_2(MatrixMuls_62_io_matA_2),
    .io_matA_3(MatrixMuls_62_io_matA_3),
    .io_matA_4(MatrixMuls_62_io_matA_4),
    .io_matA_5(MatrixMuls_62_io_matA_5),
    .io_matA_6(MatrixMuls_62_io_matA_6),
    .io_matA_7(MatrixMuls_62_io_matA_7),
    .io_matA_8(MatrixMuls_62_io_matA_8),
    .io_f_mac(MatrixMuls_62_io_f_mac)
  );
  MatMult1 MatrixMuls_63 ( // @[Convolution.scala 25:29]
    .io_matA_0(MatrixMuls_63_io_matA_0),
    .io_matA_1(MatrixMuls_63_io_matA_1),
    .io_matA_2(MatrixMuls_63_io_matA_2),
    .io_matA_3(MatrixMuls_63_io_matA_3),
    .io_matA_4(MatrixMuls_63_io_matA_4),
    .io_matA_5(MatrixMuls_63_io_matA_5),
    .io_matA_6(MatrixMuls_63_io_matA_6),
    .io_matA_7(MatrixMuls_63_io_matA_7),
    .io_matA_8(MatrixMuls_63_io_matA_8),
    .io_f_mac(MatrixMuls_63_io_f_mac)
  );
  assign io_single_out_0 = MatrixMuls_0_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_1 = MatrixMuls_1_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_2 = MatrixMuls_2_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_3 = MatrixMuls_3_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_4 = MatrixMuls_4_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_5 = MatrixMuls_5_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_6 = MatrixMuls_6_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_7 = MatrixMuls_7_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_8 = MatrixMuls_8_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_9 = MatrixMuls_9_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_10 = MatrixMuls_10_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_11 = MatrixMuls_11_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_12 = MatrixMuls_12_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_13 = MatrixMuls_13_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_14 = MatrixMuls_14_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_15 = MatrixMuls_15_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_16 = MatrixMuls_16_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_17 = MatrixMuls_17_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_18 = MatrixMuls_18_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_19 = MatrixMuls_19_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_20 = MatrixMuls_20_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_21 = MatrixMuls_21_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_22 = MatrixMuls_22_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_23 = MatrixMuls_23_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_24 = MatrixMuls_24_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_25 = MatrixMuls_25_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_26 = MatrixMuls_26_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_27 = MatrixMuls_27_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_28 = MatrixMuls_28_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_29 = MatrixMuls_29_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_30 = MatrixMuls_30_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_31 = MatrixMuls_31_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_32 = MatrixMuls_32_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_33 = MatrixMuls_33_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_34 = MatrixMuls_34_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_35 = MatrixMuls_35_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_36 = MatrixMuls_36_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_37 = MatrixMuls_37_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_38 = MatrixMuls_38_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_39 = MatrixMuls_39_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_40 = MatrixMuls_40_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_41 = MatrixMuls_41_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_42 = MatrixMuls_42_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_43 = MatrixMuls_43_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_44 = MatrixMuls_44_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_45 = MatrixMuls_45_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_46 = MatrixMuls_46_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_47 = MatrixMuls_47_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_48 = MatrixMuls_48_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_49 = MatrixMuls_49_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_50 = MatrixMuls_50_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_51 = MatrixMuls_51_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_52 = MatrixMuls_52_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_53 = MatrixMuls_53_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_54 = MatrixMuls_54_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_55 = MatrixMuls_55_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_56 = MatrixMuls_56_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_57 = MatrixMuls_57_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_58 = MatrixMuls_58_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_59 = MatrixMuls_59_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_60 = MatrixMuls_60_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_61 = MatrixMuls_61_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_62 = MatrixMuls_62_io_f_mac; // @[Convolution.scala 55:24]
  assign io_single_out_63 = MatrixMuls_63_io_f_mac; // @[Convolution.scala 55:24]
  assign MatrixMuls_0_io_matA_0 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_0_io_matA_1 = 32'h41233333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_0_io_matA_2 = 32'h4124cccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_0_io_matA_3 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_0_io_matA_4 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_0_io_matA_5 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_0_io_matA_6 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_0_io_matA_7 = 32'h404eb851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_0_io_matA_8 = 32'h410ab851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_1_io_matA_0 = 32'h41233333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_1_io_matA_1 = 32'h4124cccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_1_io_matA_2 = 32'h41266666; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_1_io_matA_3 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_1_io_matA_4 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_1_io_matA_5 = 32'h3f11eb84; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_1_io_matA_6 = 32'h404eb851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_1_io_matA_7 = 32'h410ab851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_1_io_matA_8 = 32'h411e147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_2_io_matA_0 = 32'h4124cccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_2_io_matA_1 = 32'h41266666; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_2_io_matA_2 = 32'h41280000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_2_io_matA_3 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_2_io_matA_4 = 32'h3f11eb84; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_2_io_matA_5 = 32'h3f5eb850; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_2_io_matA_6 = 32'h410ab851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_2_io_matA_7 = 32'h411e147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_2_io_matA_8 = 32'h3f47ae14; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_3_io_matA_0 = 32'h41266666; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_3_io_matA_1 = 32'h41280000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_3_io_matA_2 = 32'h41299999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_3_io_matA_3 = 32'h3f11eb84; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_3_io_matA_4 = 32'h3f5eb850; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_3_io_matA_5 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_3_io_matA_6 = 32'h411e147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_3_io_matA_7 = 32'h3f47ae14; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_3_io_matA_8 = 32'h40d147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_4_io_matA_0 = 32'h41280000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_4_io_matA_1 = 32'h41299999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_4_io_matA_2 = 32'h3ecccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_4_io_matA_3 = 32'h3f5eb850; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_4_io_matA_4 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_4_io_matA_5 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_4_io_matA_6 = 32'h3f47ae14; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_4_io_matA_7 = 32'h40d147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_4_io_matA_8 = 32'h40d80000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_5_io_matA_0 = 32'h41299999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_5_io_matA_1 = 32'h3ecccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_5_io_matA_2 = 32'h3f2e147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_5_io_matA_3 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_5_io_matA_4 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_5_io_matA_5 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_5_io_matA_6 = 32'h40d147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_5_io_matA_7 = 32'h40d80000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_5_io_matA_8 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_6_io_matA_0 = 32'h3ecccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_6_io_matA_1 = 32'h3f2e147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_6_io_matA_2 = 32'h3f6147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_6_io_matA_3 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_6_io_matA_4 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_6_io_matA_5 = 32'h3f0ccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_6_io_matA_6 = 32'h40d80000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_6_io_matA_7 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_6_io_matA_8 = 32'h40edc28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_7_io_matA_0 = 32'h3f2e147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_7_io_matA_1 = 32'h3f6147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_7_io_matA_2 = 32'h3f0ccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_7_io_matA_3 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_7_io_matA_4 = 32'h3f0ccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_7_io_matA_5 = 32'h3f9d70a3; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_7_io_matA_6 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_7_io_matA_7 = 32'h40edc28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_7_io_matA_8 = 32'h40070a3d; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_8_io_matA_0 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_8_io_matA_1 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_8_io_matA_2 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_8_io_matA_3 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_8_io_matA_4 = 32'h404eb851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_8_io_matA_5 = 32'h410ab851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_8_io_matA_6 = 32'h3f9c28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_8_io_matA_7 = 32'h3fb70a3d; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_8_io_matA_8 = 32'h40adc28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_9_io_matA_0 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_9_io_matA_1 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_9_io_matA_2 = 32'h3f11eb84; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_9_io_matA_3 = 32'h404eb851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_9_io_matA_4 = 32'h410ab851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_9_io_matA_5 = 32'h411e147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_9_io_matA_6 = 32'h3fb70a3d; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_9_io_matA_7 = 32'h40adc28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_9_io_matA_8 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_10_io_matA_0 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_10_io_matA_1 = 32'h3f11eb84; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_10_io_matA_2 = 32'h3f5eb850; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_10_io_matA_3 = 32'h410ab851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_10_io_matA_4 = 32'h411e147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_10_io_matA_5 = 32'h3f47ae14; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_10_io_matA_6 = 32'h40adc28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_10_io_matA_7 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_10_io_matA_8 = 32'h41073333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_11_io_matA_0 = 32'h3f11eb84; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_11_io_matA_1 = 32'h3f5eb850; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_11_io_matA_2 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_11_io_matA_3 = 32'h411e147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_11_io_matA_4 = 32'h3f47ae14; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_11_io_matA_5 = 32'h40d147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_11_io_matA_6 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_11_io_matA_7 = 32'h41073333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_11_io_matA_8 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_12_io_matA_0 = 32'h3f5eb850; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_12_io_matA_1 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_12_io_matA_2 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_12_io_matA_3 = 32'h3f47ae14; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_12_io_matA_4 = 32'h40d147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_12_io_matA_5 = 32'h40d80000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_12_io_matA_6 = 32'h41073333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_12_io_matA_7 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_12_io_matA_8 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_13_io_matA_0 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_13_io_matA_1 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_13_io_matA_2 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_13_io_matA_3 = 32'h40d147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_13_io_matA_4 = 32'h40d80000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_13_io_matA_5 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_13_io_matA_6 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_13_io_matA_7 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_13_io_matA_8 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_14_io_matA_0 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_14_io_matA_1 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_14_io_matA_2 = 32'h3f0ccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_14_io_matA_3 = 32'h40d80000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_14_io_matA_4 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_14_io_matA_5 = 32'h40edc28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_14_io_matA_6 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_14_io_matA_7 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_14_io_matA_8 = 32'h4114cccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_15_io_matA_0 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_15_io_matA_1 = 32'h3f0ccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_15_io_matA_2 = 32'h3f9d70a3; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_15_io_matA_3 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_15_io_matA_4 = 32'h40edc28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_15_io_matA_5 = 32'h40070a3d; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_15_io_matA_6 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_15_io_matA_7 = 32'h4114cccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_15_io_matA_8 = 32'h3fb33333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_16_io_matA_0 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_16_io_matA_1 = 32'h404eb851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_16_io_matA_2 = 32'h410ab851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_16_io_matA_3 = 32'h3f9c28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_16_io_matA_4 = 32'h3fb70a3d; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_16_io_matA_5 = 32'h40adc28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_16_io_matA_6 = 32'h3fc00000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_16_io_matA_7 = 32'h40266666; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_16_io_matA_8 = 32'h40599999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_17_io_matA_0 = 32'h404eb851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_17_io_matA_1 = 32'h410ab851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_17_io_matA_2 = 32'h411e147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_17_io_matA_3 = 32'h3fb70a3d; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_17_io_matA_4 = 32'h40adc28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_17_io_matA_5 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_17_io_matA_6 = 32'h40266666; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_17_io_matA_7 = 32'h40599999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_17_io_matA_8 = 32'h40b5c28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_18_io_matA_0 = 32'h410ab851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_18_io_matA_1 = 32'h411e147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_18_io_matA_2 = 32'h3f47ae14; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_18_io_matA_3 = 32'h40adc28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_18_io_matA_4 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_18_io_matA_5 = 32'h41073333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_18_io_matA_6 = 32'h40599999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_18_io_matA_7 = 32'h40b5c28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_18_io_matA_8 = 32'h40fc28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_19_io_matA_0 = 32'h411e147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_19_io_matA_1 = 32'h3f47ae14; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_19_io_matA_2 = 32'h40d147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_19_io_matA_3 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_19_io_matA_4 = 32'h41073333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_19_io_matA_5 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_19_io_matA_6 = 32'h40b5c28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_19_io_matA_7 = 32'h40fc28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_19_io_matA_8 = 32'h40919999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_20_io_matA_0 = 32'h3f47ae14; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_20_io_matA_1 = 32'h40d147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_20_io_matA_2 = 32'h40d80000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_20_io_matA_3 = 32'h41073333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_20_io_matA_4 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_20_io_matA_5 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_20_io_matA_6 = 32'h40fc28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_20_io_matA_7 = 32'h40919999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_20_io_matA_8 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_21_io_matA_0 = 32'h40d147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_21_io_matA_1 = 32'h40d80000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_21_io_matA_2 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_21_io_matA_3 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_21_io_matA_4 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_21_io_matA_5 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_21_io_matA_6 = 32'h40919999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_21_io_matA_7 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_21_io_matA_8 = 32'h401c28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_22_io_matA_0 = 32'h40d80000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_22_io_matA_1 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_22_io_matA_2 = 32'h40edc28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_22_io_matA_3 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_22_io_matA_4 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_22_io_matA_5 = 32'h4114cccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_22_io_matA_6 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_22_io_matA_7 = 32'h401c28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_22_io_matA_8 = 32'h40ae147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_23_io_matA_0 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_23_io_matA_1 = 32'h40edc28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_23_io_matA_2 = 32'h40070a3d; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_23_io_matA_3 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_23_io_matA_4 = 32'h4114cccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_23_io_matA_5 = 32'h3fb33333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_23_io_matA_6 = 32'h401c28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_23_io_matA_7 = 32'h40ae147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_23_io_matA_8 = 32'h40d23d70; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_24_io_matA_0 = 32'h3f9c28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_24_io_matA_1 = 32'h3fb70a3d; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_24_io_matA_2 = 32'h40adc28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_24_io_matA_3 = 32'h3fc00000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_24_io_matA_4 = 32'h40266666; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_24_io_matA_5 = 32'h40599999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_24_io_matA_6 = 32'h410deb85; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_24_io_matA_7 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_24_io_matA_8 = 32'h40551eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_25_io_matA_0 = 32'h3fb70a3d; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_25_io_matA_1 = 32'h40adc28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_25_io_matA_2 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_25_io_matA_3 = 32'h40266666; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_25_io_matA_4 = 32'h40599999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_25_io_matA_5 = 32'h40b5c28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_25_io_matA_6 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_25_io_matA_7 = 32'h40551eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_25_io_matA_8 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_26_io_matA_0 = 32'h40adc28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_26_io_matA_1 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_26_io_matA_2 = 32'h41073333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_26_io_matA_3 = 32'h40599999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_26_io_matA_4 = 32'h40b5c28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_26_io_matA_5 = 32'h40fc28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_26_io_matA_6 = 32'h40551eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_26_io_matA_7 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_26_io_matA_8 = 32'h40b19999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_27_io_matA_0 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_27_io_matA_1 = 32'h41073333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_27_io_matA_2 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_27_io_matA_3 = 32'h40b5c28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_27_io_matA_4 = 32'h40fc28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_27_io_matA_5 = 32'h40919999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_27_io_matA_6 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_27_io_matA_7 = 32'h40b19999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_27_io_matA_8 = 32'h3f9d70a3; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_28_io_matA_0 = 32'h41073333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_28_io_matA_1 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_28_io_matA_2 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_28_io_matA_3 = 32'h40fc28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_28_io_matA_4 = 32'h40919999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_28_io_matA_5 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_28_io_matA_6 = 32'h40b19999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_28_io_matA_7 = 32'h3f9d70a3; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_28_io_matA_8 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_29_io_matA_0 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_29_io_matA_1 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_29_io_matA_2 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_29_io_matA_3 = 32'h40919999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_29_io_matA_4 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_29_io_matA_5 = 32'h401c28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_29_io_matA_6 = 32'h3f9d70a3; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_29_io_matA_7 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_29_io_matA_8 = 32'h404eb851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_30_io_matA_0 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_30_io_matA_1 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_30_io_matA_2 = 32'h4114cccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_30_io_matA_3 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_30_io_matA_4 = 32'h401c28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_30_io_matA_5 = 32'h40ae147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_30_io_matA_6 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_30_io_matA_7 = 32'h404eb851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_30_io_matA_8 = 32'h3f2b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_31_io_matA_0 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_31_io_matA_1 = 32'h4114cccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_31_io_matA_2 = 32'h3fb33333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_31_io_matA_3 = 32'h401c28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_31_io_matA_4 = 32'h40ae147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_31_io_matA_5 = 32'h40d23d70; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_31_io_matA_6 = 32'h404eb851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_31_io_matA_7 = 32'h3f2b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_31_io_matA_8 = 32'h3f6147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_32_io_matA_0 = 32'h3fc00000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_32_io_matA_1 = 32'h40266666; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_32_io_matA_2 = 32'h40599999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_32_io_matA_3 = 32'h410deb85; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_32_io_matA_4 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_32_io_matA_5 = 32'h40551eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_32_io_matA_6 = 32'h3f47ae14; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_32_io_matA_7 = 32'h3f0a3d70; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_32_io_matA_8 = 32'h3f400000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_33_io_matA_0 = 32'h40266666; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_33_io_matA_1 = 32'h40599999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_33_io_matA_2 = 32'h40b5c28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_33_io_matA_3 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_33_io_matA_4 = 32'h40551eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_33_io_matA_5 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_33_io_matA_6 = 32'h3f0a3d70; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_33_io_matA_7 = 32'h3f400000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_33_io_matA_8 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_34_io_matA_0 = 32'h40599999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_34_io_matA_1 = 32'h40b5c28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_34_io_matA_2 = 32'h40fc28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_34_io_matA_3 = 32'h40551eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_34_io_matA_4 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_34_io_matA_5 = 32'h40b19999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_34_io_matA_6 = 32'h3f400000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_34_io_matA_7 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_34_io_matA_8 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_35_io_matA_0 = 32'h40b5c28f; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_35_io_matA_1 = 32'h40fc28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_35_io_matA_2 = 32'h40919999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_35_io_matA_3 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_35_io_matA_4 = 32'h40b19999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_35_io_matA_5 = 32'h3f9d70a3; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_35_io_matA_6 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_35_io_matA_7 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_35_io_matA_8 = 32'h3de147a0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_36_io_matA_0 = 32'h40fc28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_36_io_matA_1 = 32'h40919999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_36_io_matA_2 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_36_io_matA_3 = 32'h40b19999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_36_io_matA_4 = 32'h3f9d70a3; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_36_io_matA_5 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_36_io_matA_6 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_36_io_matA_7 = 32'h3de147a0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_36_io_matA_8 = 32'h3e6147a8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_37_io_matA_0 = 32'h40919999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_37_io_matA_1 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_37_io_matA_2 = 32'h401c28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_37_io_matA_3 = 32'h3f9d70a3; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_37_io_matA_4 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_37_io_matA_5 = 32'h404eb851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_37_io_matA_6 = 32'h3de147a0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_37_io_matA_7 = 32'h3e6147a8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_37_io_matA_8 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_38_io_matA_0 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_38_io_matA_1 = 32'h401c28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_38_io_matA_2 = 32'h40ae147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_38_io_matA_3 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_38_io_matA_4 = 32'h404eb851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_38_io_matA_5 = 32'h3f2b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_38_io_matA_6 = 32'h3e6147a8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_38_io_matA_7 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_38_io_matA_8 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_39_io_matA_0 = 32'h401c28f5; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_39_io_matA_1 = 32'h40ae147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_39_io_matA_2 = 32'h40d23d70; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_39_io_matA_3 = 32'h404eb851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_39_io_matA_4 = 32'h3f2b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_39_io_matA_5 = 32'h3f6147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_39_io_matA_6 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_39_io_matA_7 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_39_io_matA_8 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_40_io_matA_0 = 32'h410deb85; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_40_io_matA_1 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_40_io_matA_2 = 32'h40551eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_40_io_matA_3 = 32'h3f47ae14; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_40_io_matA_4 = 32'h3f0a3d70; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_40_io_matA_5 = 32'h3f400000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_40_io_matA_6 = 32'h3ee66664; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_40_io_matA_7 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_40_io_matA_8 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_41_io_matA_0 = 32'h40d8a3d7; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_41_io_matA_1 = 32'h40551eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_41_io_matA_2 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_41_io_matA_3 = 32'h3f0a3d70; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_41_io_matA_4 = 32'h3f400000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_41_io_matA_5 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_41_io_matA_6 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_41_io_matA_7 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_41_io_matA_8 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_42_io_matA_0 = 32'h40551eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_42_io_matA_1 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_42_io_matA_2 = 32'h40b19999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_42_io_matA_3 = 32'h3f400000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_42_io_matA_4 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_42_io_matA_5 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_42_io_matA_6 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_42_io_matA_7 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_42_io_matA_8 = 32'h3e999998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_43_io_matA_0 = 32'h40151eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_43_io_matA_1 = 32'h40b19999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_43_io_matA_2 = 32'h3f9d70a3; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_43_io_matA_3 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_43_io_matA_4 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_43_io_matA_5 = 32'h3de147a0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_43_io_matA_6 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_43_io_matA_7 = 32'h3e999998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_43_io_matA_8 = 32'h3fb33333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_44_io_matA_0 = 32'h40b19999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_44_io_matA_1 = 32'h3f9d70a3; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_44_io_matA_2 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_44_io_matA_3 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_44_io_matA_4 = 32'h3de147a0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_44_io_matA_5 = 32'h3e6147a8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_44_io_matA_6 = 32'h3e999998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_44_io_matA_7 = 32'h3fb33333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_44_io_matA_8 = 32'h3f000000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_45_io_matA_0 = 32'h3f9d70a3; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_45_io_matA_1 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_45_io_matA_2 = 32'h404eb851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_45_io_matA_3 = 32'h3de147a0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_45_io_matA_4 = 32'h3e6147a8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_45_io_matA_5 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_45_io_matA_6 = 32'h3fb33333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_45_io_matA_7 = 32'h3f000000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_45_io_matA_8 = 32'h3f199998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_46_io_matA_0 = 32'h405b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_46_io_matA_1 = 32'h404eb851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_46_io_matA_2 = 32'h3f2b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_46_io_matA_3 = 32'h3e6147a8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_46_io_matA_4 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_46_io_matA_5 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_46_io_matA_6 = 32'h3f000000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_46_io_matA_7 = 32'h3f199998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_46_io_matA_8 = 32'h3ecccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_47_io_matA_0 = 32'h404eb851; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_47_io_matA_1 = 32'h3f2b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_47_io_matA_2 = 32'h3f6147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_47_io_matA_3 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_47_io_matA_4 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_47_io_matA_5 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_47_io_matA_6 = 32'h3f199998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_47_io_matA_7 = 32'h3ecccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_47_io_matA_8 = 32'h3f2e147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_48_io_matA_0 = 32'h3f47ae14; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_48_io_matA_1 = 32'h3f0a3d70; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_48_io_matA_2 = 32'h3f400000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_48_io_matA_3 = 32'h3ee66664; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_48_io_matA_4 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_48_io_matA_5 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_48_io_matA_6 = 32'h3f6147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_48_io_matA_7 = 32'h3f0ccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_48_io_matA_8 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_49_io_matA_0 = 32'h3f0a3d70; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_49_io_matA_1 = 32'h3f400000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_49_io_matA_2 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_49_io_matA_3 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_49_io_matA_4 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_49_io_matA_5 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_49_io_matA_6 = 32'h3f0ccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_49_io_matA_7 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_49_io_matA_8 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_50_io_matA_0 = 32'h3f400000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_50_io_matA_1 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_50_io_matA_2 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_50_io_matA_3 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_50_io_matA_4 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_50_io_matA_5 = 32'h3e999998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_50_io_matA_6 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_50_io_matA_7 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_50_io_matA_8 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_51_io_matA_0 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_51_io_matA_1 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_51_io_matA_2 = 32'h3de147a0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_51_io_matA_3 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_51_io_matA_4 = 32'h3e999998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_51_io_matA_5 = 32'h3fb33333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_51_io_matA_6 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_51_io_matA_7 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_51_io_matA_8 = 32'h3f11eb84; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_52_io_matA_0 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_52_io_matA_1 = 32'h3de147a0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_52_io_matA_2 = 32'h3e6147a8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_52_io_matA_3 = 32'h3e999998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_52_io_matA_4 = 32'h3fb33333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_52_io_matA_5 = 32'h3f000000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_52_io_matA_6 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_52_io_matA_7 = 32'h3f11eb84; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_52_io_matA_8 = 32'h3f5eb850; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_53_io_matA_0 = 32'h3de147a0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_53_io_matA_1 = 32'h3e6147a8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_53_io_matA_2 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_53_io_matA_3 = 32'h3fb33333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_53_io_matA_4 = 32'h3f000000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_53_io_matA_5 = 32'h3f199998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_53_io_matA_6 = 32'h3f11eb84; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_53_io_matA_7 = 32'h3f5eb850; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_53_io_matA_8 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_54_io_matA_0 = 32'h3e6147a8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_54_io_matA_1 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_54_io_matA_2 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_54_io_matA_3 = 32'h3f000000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_54_io_matA_4 = 32'h3f199998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_54_io_matA_5 = 32'h3ecccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_54_io_matA_6 = 32'h3f5eb850; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_54_io_matA_7 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_54_io_matA_8 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_55_io_matA_0 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_55_io_matA_1 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_55_io_matA_2 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_55_io_matA_3 = 32'h3f199998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_55_io_matA_4 = 32'h3ecccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_55_io_matA_5 = 32'h3f2e147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_55_io_matA_6 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_55_io_matA_7 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_55_io_matA_8 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_56_io_matA_0 = 32'h3ee66664; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_56_io_matA_1 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_56_io_matA_2 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_56_io_matA_3 = 32'h3f6147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_56_io_matA_4 = 32'h3f0ccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_56_io_matA_5 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_56_io_matA_6 = 32'h3f0ccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_56_io_matA_7 = 32'h3e6b8518; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_56_io_matA_8 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_57_io_matA_0 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_57_io_matA_1 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_57_io_matA_2 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_57_io_matA_3 = 32'h3f0ccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_57_io_matA_4 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_57_io_matA_5 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_57_io_matA_6 = 32'h3e6b8518; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_57_io_matA_7 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_57_io_matA_8 = 32'h3e6b8518; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_58_io_matA_0 = 32'h3dccccc0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_58_io_matA_1 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_58_io_matA_2 = 32'h3e999998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_58_io_matA_3 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_58_io_matA_4 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_58_io_matA_5 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_58_io_matA_6 = 32'h3edc28f4; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_58_io_matA_7 = 32'h3e6b8518; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_58_io_matA_8 = 32'h3f2b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_59_io_matA_0 = 32'h3f999999; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_59_io_matA_1 = 32'h3e999998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_59_io_matA_2 = 32'h3fb33333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_59_io_matA_3 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_59_io_matA_4 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_59_io_matA_5 = 32'h3f11eb84; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_59_io_matA_6 = 32'h3e6b8518; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_59_io_matA_7 = 32'h3f2b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_59_io_matA_8 = 32'h3f6147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_60_io_matA_0 = 32'h3e999998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_60_io_matA_1 = 32'h3fb33333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_60_io_matA_2 = 32'h3f000000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_60_io_matA_3 = 32'h3ee147ac; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_60_io_matA_4 = 32'h3f11eb84; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_60_io_matA_5 = 32'h3f5eb850; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_60_io_matA_6 = 32'h3f2b851e; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_60_io_matA_7 = 32'h3f6147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_60_io_matA_8 = 32'h3f47ae14; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_61_io_matA_0 = 32'h3fb33333; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_61_io_matA_1 = 32'h3f000000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_61_io_matA_2 = 32'h3f199998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_61_io_matA_3 = 32'h3f11eb84; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_61_io_matA_4 = 32'h3f5eb850; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_61_io_matA_5 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_61_io_matA_6 = 32'h3f6147ae; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_61_io_matA_7 = 32'h3f47ae14; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_61_io_matA_8 = 32'h3f0a3d70; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_62_io_matA_0 = 32'h3f000000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_62_io_matA_1 = 32'h3f199998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_62_io_matA_2 = 32'h3ecccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_62_io_matA_3 = 32'h3f5eb850; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_62_io_matA_4 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_62_io_matA_5 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_62_io_matA_6 = 32'h3f47ae14; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_62_io_matA_7 = 32'h3f0a3d70; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_62_io_matA_8 = 32'h3f400000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_63_io_matA_0 = 32'h3f199998; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_63_io_matA_1 = 32'h3ecccccc; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_63_io_matA_2 = 32'h3f2e147a; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_63_io_matA_3 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_63_io_matA_4 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_63_io_matA_5 = 32'h3ea8f5c0; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_63_io_matA_6 = 32'h3f0a3d70; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_63_io_matA_7 = 32'h3f400000; // @[Convolution.scala 35:22 43:27]
  assign MatrixMuls_63_io_matA_8 = 32'h3f451eb8; // @[Convolution.scala 35:22 43:27]
endmodule
module full_subber_1729(
  input  [22:0] io_in_a,
  input  [22:0] io_in_b,
  output        io_out_c
);
  wire [23:0] _result_T = io_in_a - io_in_b; // @[Arithmetic.scala 70:23]
  wire [24:0] _result_T_2 = _result_T - 24'h0; // @[Arithmetic.scala 70:34]
  wire [23:0] result = _result_T_2[23:0]; // @[Arithmetic.scala 69:22 70:12]
  assign io_out_c = result[23]; // @[Arithmetic.scala 72:23]
endmodule
module FP_Comparitor(
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
  wire [7:0] full_subber_io_in_a; // @[FPArithmetic.scala 777:24]
  wire [7:0] full_subber_io_in_b; // @[FPArithmetic.scala 777:24]
  wire [7:0] full_subber_io_out_s; // @[FPArithmetic.scala 777:24]
  wire  full_subber_io_out_c; // @[FPArithmetic.scala 777:24]
  wire [22:0] full_subber_1_io_in_a; // @[FPArithmetic.scala 782:25]
  wire [22:0] full_subber_1_io_in_b; // @[FPArithmetic.scala 782:25]
  wire  full_subber_1_io_out_c; // @[FPArithmetic.scala 782:25]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FPArithmetic.scala 756:62]
  wire [8:0] _GEN_5 = {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 756:34]
  wire [8:0] _GEN_0 = _GEN_5 > _T_2 ? _T_2 : {{1'd0}, io_in_a[30:23]}; // @[FPArithmetic.scala 756:68 757:14 759:14]
  wire [8:0] _GEN_6 = {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 761:34]
  wire [8:0] _GEN_1 = _GEN_6 > _T_2 ? _T_2 : {{1'd0}, io_in_b[30:23]}; // @[FPArithmetic.scala 761:68 762:14 764:14]
  wire [31:0] _GEN_2 = full_subber_1_io_out_c ? io_in_b : io_in_a; // @[FPArithmetic.scala 792:34 793:18 795:18]
  wire [31:0] _GEN_3 = full_subber_io_out_s > 8'h0 ? io_in_a : _GEN_2; // @[FPArithmetic.scala 789:35 790:16]
  full_subber full_subber ( // @[FPArithmetic.scala 777:24]
    .io_in_a(full_subber_io_in_a),
    .io_in_b(full_subber_io_in_b),
    .io_out_s(full_subber_io_out_s),
    .io_out_c(full_subber_io_out_c)
  );
  full_subber_1729 full_subber_1 ( // @[FPArithmetic.scala 782:25]
    .io_in_a(full_subber_1_io_in_a),
    .io_in_b(full_subber_1_io_in_b),
    .io_out_c(full_subber_1_io_out_c)
  );
  assign io_out_s = full_subber_io_out_c ? io_in_b : _GEN_3; // @[FPArithmetic.scala 787:31 788:16]
  assign full_subber_io_in_a = _GEN_0[7:0]; // @[FPArithmetic.scala 755:19]
  assign full_subber_io_in_b = _GEN_1[7:0]; // @[FPArithmetic.scala 755:19]
  assign full_subber_1_io_in_a = io_in_a[22:0]; // @[FPArithmetic.scala 769:23]
  assign full_subber_1_io_in_b = io_in_b[22:0]; // @[FPArithmetic.scala 770:23]
endmodule
module Max_Pooling(
  input  [31:0] io_pixel1,
  input  [31:0] io_pixel2,
  input  [31:0] io_pixel3,
  input  [31:0] io_pixel4,
  output [31:0] io_f_max
);
  wire [31:0] fp1_io_in_a; // @[Pooling.scala 19:21]
  wire [31:0] fp1_io_in_b; // @[Pooling.scala 19:21]
  wire [31:0] fp1_io_out_s; // @[Pooling.scala 19:21]
  wire [31:0] fp2_io_in_a; // @[Pooling.scala 24:21]
  wire [31:0] fp2_io_in_b; // @[Pooling.scala 24:21]
  wire [31:0] fp2_io_out_s; // @[Pooling.scala 24:21]
  wire [31:0] fp3_io_in_a; // @[Pooling.scala 29:21]
  wire [31:0] fp3_io_in_b; // @[Pooling.scala 29:21]
  wire [31:0] fp3_io_out_s; // @[Pooling.scala 29:21]
  FP_Comparitor fp1 ( // @[Pooling.scala 19:21]
    .io_in_a(fp1_io_in_a),
    .io_in_b(fp1_io_in_b),
    .io_out_s(fp1_io_out_s)
  );
  FP_Comparitor fp2 ( // @[Pooling.scala 24:21]
    .io_in_a(fp2_io_in_a),
    .io_in_b(fp2_io_in_b),
    .io_out_s(fp2_io_out_s)
  );
  FP_Comparitor fp3 ( // @[Pooling.scala 29:21]
    .io_in_a(fp3_io_in_a),
    .io_in_b(fp3_io_in_b),
    .io_out_s(fp3_io_out_s)
  );
  assign io_f_max = fp3_io_out_s; // @[Pooling.scala 32:14]
  assign fp1_io_in_a = io_pixel1; // @[Pooling.scala 20:17]
  assign fp1_io_in_b = io_pixel2; // @[Pooling.scala 21:17]
  assign fp2_io_in_a = io_pixel3; // @[Pooling.scala 25:17]
  assign fp2_io_in_b = io_pixel4; // @[Pooling.scala 26:17]
  assign fp3_io_in_a = fp1_io_out_s; // @[Pooling.scala 16:20 22:10]
  assign fp3_io_in_b = fp2_io_out_s; // @[Pooling.scala 17:20 27:10]
endmodule
module Pooling_Controller(
  input         clock,
  input  [31:0] io_InputMatrix_0,
  input  [31:0] io_InputMatrix_1,
  input  [31:0] io_InputMatrix_2,
  input  [31:0] io_InputMatrix_3,
  input  [31:0] io_InputMatrix_4,
  input  [31:0] io_InputMatrix_5,
  input  [31:0] io_InputMatrix_6,
  input  [31:0] io_InputMatrix_7,
  input  [31:0] io_InputMatrix_8,
  input  [31:0] io_InputMatrix_9,
  input  [31:0] io_InputMatrix_10,
  input  [31:0] io_InputMatrix_11,
  input  [31:0] io_InputMatrix_12,
  input  [31:0] io_InputMatrix_13,
  input  [31:0] io_InputMatrix_14,
  input  [31:0] io_InputMatrix_15,
  input  [31:0] io_InputMatrix_16,
  input  [31:0] io_InputMatrix_17,
  input  [31:0] io_InputMatrix_18,
  input  [31:0] io_InputMatrix_19,
  input  [31:0] io_InputMatrix_20,
  input  [31:0] io_InputMatrix_21,
  input  [31:0] io_InputMatrix_22,
  input  [31:0] io_InputMatrix_23,
  input  [31:0] io_InputMatrix_24,
  input  [31:0] io_InputMatrix_25,
  input  [31:0] io_InputMatrix_26,
  input  [31:0] io_InputMatrix_27,
  input  [31:0] io_InputMatrix_28,
  input  [31:0] io_InputMatrix_29,
  input  [31:0] io_InputMatrix_30,
  input  [31:0] io_InputMatrix_31,
  input  [31:0] io_InputMatrix_32,
  input  [31:0] io_InputMatrix_33,
  input  [31:0] io_InputMatrix_34,
  input  [31:0] io_InputMatrix_35,
  input  [31:0] io_InputMatrix_36,
  input  [31:0] io_InputMatrix_37,
  input  [31:0] io_InputMatrix_38,
  input  [31:0] io_InputMatrix_39,
  input  [31:0] io_InputMatrix_40,
  input  [31:0] io_InputMatrix_41,
  input  [31:0] io_InputMatrix_42,
  input  [31:0] io_InputMatrix_43,
  input  [31:0] io_InputMatrix_44,
  input  [31:0] io_InputMatrix_45,
  input  [31:0] io_InputMatrix_46,
  input  [31:0] io_InputMatrix_47,
  input  [31:0] io_InputMatrix_48,
  input  [31:0] io_InputMatrix_49,
  input  [31:0] io_InputMatrix_50,
  input  [31:0] io_InputMatrix_51,
  input  [31:0] io_InputMatrix_52,
  input  [31:0] io_InputMatrix_53,
  input  [31:0] io_InputMatrix_54,
  input  [31:0] io_InputMatrix_55,
  input  [31:0] io_InputMatrix_56,
  input  [31:0] io_InputMatrix_57,
  input  [31:0] io_InputMatrix_58,
  input  [31:0] io_InputMatrix_59,
  input  [31:0] io_InputMatrix_60,
  input  [31:0] io_InputMatrix_61,
  input  [31:0] io_InputMatrix_62,
  input  [31:0] io_InputMatrix_63,
  output [31:0] io_single_out_0,
  output [31:0] io_single_out_1,
  output [31:0] io_single_out_2,
  output [31:0] io_single_out_3,
  output [31:0] io_single_out_4,
  output [31:0] io_single_out_5,
  output [31:0] io_single_out_6,
  output [31:0] io_single_out_7,
  output [31:0] io_single_out_8,
  output [31:0] io_single_out_9,
  output [31:0] io_single_out_10,
  output [31:0] io_single_out_11,
  output [31:0] io_single_out_12,
  output [31:0] io_single_out_13,
  output [31:0] io_single_out_14,
  output [31:0] io_single_out_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] Max_Poolings_0_io_pixel1; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_0_io_pixel2; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_0_io_pixel3; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_0_io_pixel4; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_0_io_f_max; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_1_io_pixel1; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_1_io_pixel2; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_1_io_pixel3; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_1_io_pixel4; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_1_io_f_max; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_2_io_pixel1; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_2_io_pixel2; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_2_io_pixel3; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_2_io_pixel4; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_2_io_f_max; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_3_io_pixel1; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_3_io_pixel2; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_3_io_pixel3; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_3_io_pixel4; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_3_io_f_max; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_4_io_pixel1; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_4_io_pixel2; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_4_io_pixel3; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_4_io_pixel4; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_4_io_f_max; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_5_io_pixel1; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_5_io_pixel2; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_5_io_pixel3; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_5_io_pixel4; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_5_io_f_max; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_6_io_pixel1; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_6_io_pixel2; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_6_io_pixel3; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_6_io_pixel4; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_6_io_f_max; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_7_io_pixel1; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_7_io_pixel2; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_7_io_pixel3; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_7_io_pixel4; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_7_io_f_max; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_8_io_pixel1; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_8_io_pixel2; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_8_io_pixel3; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_8_io_pixel4; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_8_io_f_max; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_9_io_pixel1; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_9_io_pixel2; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_9_io_pixel3; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_9_io_pixel4; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_9_io_f_max; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_10_io_pixel1; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_10_io_pixel2; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_10_io_pixel3; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_10_io_pixel4; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_10_io_f_max; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_11_io_pixel1; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_11_io_pixel2; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_11_io_pixel3; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_11_io_pixel4; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_11_io_f_max; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_12_io_pixel1; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_12_io_pixel2; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_12_io_pixel3; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_12_io_pixel4; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_12_io_f_max; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_13_io_pixel1; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_13_io_pixel2; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_13_io_pixel3; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_13_io_pixel4; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_13_io_f_max; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_14_io_pixel1; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_14_io_pixel2; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_14_io_pixel3; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_14_io_pixel4; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_14_io_f_max; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_15_io_pixel1; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_15_io_pixel2; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_15_io_pixel3; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_15_io_pixel4; // @[PoolingController.scala 23:31]
  wire [31:0] Max_Poolings_15_io_f_max; // @[PoolingController.scala 23:31]
  reg [31:0] values_0; // @[PoolingController.scala 20:21]
  reg [31:0] values_1; // @[PoolingController.scala 20:21]
  reg [31:0] values_2; // @[PoolingController.scala 20:21]
  reg [31:0] values_3; // @[PoolingController.scala 20:21]
  reg [31:0] values_4; // @[PoolingController.scala 20:21]
  reg [31:0] values_5; // @[PoolingController.scala 20:21]
  reg [31:0] values_6; // @[PoolingController.scala 20:21]
  reg [31:0] values_7; // @[PoolingController.scala 20:21]
  reg [31:0] values_8; // @[PoolingController.scala 20:21]
  reg [31:0] values_9; // @[PoolingController.scala 20:21]
  reg [31:0] values_10; // @[PoolingController.scala 20:21]
  reg [31:0] values_11; // @[PoolingController.scala 20:21]
  reg [31:0] values_12; // @[PoolingController.scala 20:21]
  reg [31:0] values_13; // @[PoolingController.scala 20:21]
  reg [31:0] values_14; // @[PoolingController.scala 20:21]
  reg [31:0] values_15; // @[PoolingController.scala 20:21]
  reg [31:0] values_16; // @[PoolingController.scala 20:21]
  reg [31:0] values_17; // @[PoolingController.scala 20:21]
  reg [31:0] values_18; // @[PoolingController.scala 20:21]
  reg [31:0] values_19; // @[PoolingController.scala 20:21]
  reg [31:0] values_20; // @[PoolingController.scala 20:21]
  reg [31:0] values_21; // @[PoolingController.scala 20:21]
  reg [31:0] values_22; // @[PoolingController.scala 20:21]
  reg [31:0] values_23; // @[PoolingController.scala 20:21]
  reg [31:0] values_24; // @[PoolingController.scala 20:21]
  reg [31:0] values_25; // @[PoolingController.scala 20:21]
  reg [31:0] values_26; // @[PoolingController.scala 20:21]
  reg [31:0] values_27; // @[PoolingController.scala 20:21]
  reg [31:0] values_28; // @[PoolingController.scala 20:21]
  reg [31:0] values_29; // @[PoolingController.scala 20:21]
  reg [31:0] values_30; // @[PoolingController.scala 20:21]
  reg [31:0] values_31; // @[PoolingController.scala 20:21]
  reg [31:0] values_32; // @[PoolingController.scala 20:21]
  reg [31:0] values_33; // @[PoolingController.scala 20:21]
  reg [31:0] values_34; // @[PoolingController.scala 20:21]
  reg [31:0] values_35; // @[PoolingController.scala 20:21]
  reg [31:0] values_36; // @[PoolingController.scala 20:21]
  reg [31:0] values_37; // @[PoolingController.scala 20:21]
  reg [31:0] values_38; // @[PoolingController.scala 20:21]
  reg [31:0] values_39; // @[PoolingController.scala 20:21]
  reg [31:0] values_40; // @[PoolingController.scala 20:21]
  reg [31:0] values_41; // @[PoolingController.scala 20:21]
  reg [31:0] values_42; // @[PoolingController.scala 20:21]
  reg [31:0] values_43; // @[PoolingController.scala 20:21]
  reg [31:0] values_44; // @[PoolingController.scala 20:21]
  reg [31:0] values_45; // @[PoolingController.scala 20:21]
  reg [31:0] values_46; // @[PoolingController.scala 20:21]
  reg [31:0] values_47; // @[PoolingController.scala 20:21]
  reg [31:0] values_48; // @[PoolingController.scala 20:21]
  reg [31:0] values_49; // @[PoolingController.scala 20:21]
  reg [31:0] values_50; // @[PoolingController.scala 20:21]
  reg [31:0] values_51; // @[PoolingController.scala 20:21]
  reg [31:0] values_52; // @[PoolingController.scala 20:21]
  reg [31:0] values_53; // @[PoolingController.scala 20:21]
  reg [31:0] values_54; // @[PoolingController.scala 20:21]
  reg [31:0] values_55; // @[PoolingController.scala 20:21]
  reg [31:0] values_56; // @[PoolingController.scala 20:21]
  reg [31:0] values_57; // @[PoolingController.scala 20:21]
  reg [31:0] values_58; // @[PoolingController.scala 20:21]
  reg [31:0] values_59; // @[PoolingController.scala 20:21]
  reg [31:0] values_60; // @[PoolingController.scala 20:21]
  reg [31:0] values_61; // @[PoolingController.scala 20:21]
  reg [31:0] values_62; // @[PoolingController.scala 20:21]
  reg [31:0] values_63; // @[PoolingController.scala 20:21]
  Max_Pooling Max_Poolings_0 ( // @[PoolingController.scala 23:31]
    .io_pixel1(Max_Poolings_0_io_pixel1),
    .io_pixel2(Max_Poolings_0_io_pixel2),
    .io_pixel3(Max_Poolings_0_io_pixel3),
    .io_pixel4(Max_Poolings_0_io_pixel4),
    .io_f_max(Max_Poolings_0_io_f_max)
  );
  Max_Pooling Max_Poolings_1 ( // @[PoolingController.scala 23:31]
    .io_pixel1(Max_Poolings_1_io_pixel1),
    .io_pixel2(Max_Poolings_1_io_pixel2),
    .io_pixel3(Max_Poolings_1_io_pixel3),
    .io_pixel4(Max_Poolings_1_io_pixel4),
    .io_f_max(Max_Poolings_1_io_f_max)
  );
  Max_Pooling Max_Poolings_2 ( // @[PoolingController.scala 23:31]
    .io_pixel1(Max_Poolings_2_io_pixel1),
    .io_pixel2(Max_Poolings_2_io_pixel2),
    .io_pixel3(Max_Poolings_2_io_pixel3),
    .io_pixel4(Max_Poolings_2_io_pixel4),
    .io_f_max(Max_Poolings_2_io_f_max)
  );
  Max_Pooling Max_Poolings_3 ( // @[PoolingController.scala 23:31]
    .io_pixel1(Max_Poolings_3_io_pixel1),
    .io_pixel2(Max_Poolings_3_io_pixel2),
    .io_pixel3(Max_Poolings_3_io_pixel3),
    .io_pixel4(Max_Poolings_3_io_pixel4),
    .io_f_max(Max_Poolings_3_io_f_max)
  );
  Max_Pooling Max_Poolings_4 ( // @[PoolingController.scala 23:31]
    .io_pixel1(Max_Poolings_4_io_pixel1),
    .io_pixel2(Max_Poolings_4_io_pixel2),
    .io_pixel3(Max_Poolings_4_io_pixel3),
    .io_pixel4(Max_Poolings_4_io_pixel4),
    .io_f_max(Max_Poolings_4_io_f_max)
  );
  Max_Pooling Max_Poolings_5 ( // @[PoolingController.scala 23:31]
    .io_pixel1(Max_Poolings_5_io_pixel1),
    .io_pixel2(Max_Poolings_5_io_pixel2),
    .io_pixel3(Max_Poolings_5_io_pixel3),
    .io_pixel4(Max_Poolings_5_io_pixel4),
    .io_f_max(Max_Poolings_5_io_f_max)
  );
  Max_Pooling Max_Poolings_6 ( // @[PoolingController.scala 23:31]
    .io_pixel1(Max_Poolings_6_io_pixel1),
    .io_pixel2(Max_Poolings_6_io_pixel2),
    .io_pixel3(Max_Poolings_6_io_pixel3),
    .io_pixel4(Max_Poolings_6_io_pixel4),
    .io_f_max(Max_Poolings_6_io_f_max)
  );
  Max_Pooling Max_Poolings_7 ( // @[PoolingController.scala 23:31]
    .io_pixel1(Max_Poolings_7_io_pixel1),
    .io_pixel2(Max_Poolings_7_io_pixel2),
    .io_pixel3(Max_Poolings_7_io_pixel3),
    .io_pixel4(Max_Poolings_7_io_pixel4),
    .io_f_max(Max_Poolings_7_io_f_max)
  );
  Max_Pooling Max_Poolings_8 ( // @[PoolingController.scala 23:31]
    .io_pixel1(Max_Poolings_8_io_pixel1),
    .io_pixel2(Max_Poolings_8_io_pixel2),
    .io_pixel3(Max_Poolings_8_io_pixel3),
    .io_pixel4(Max_Poolings_8_io_pixel4),
    .io_f_max(Max_Poolings_8_io_f_max)
  );
  Max_Pooling Max_Poolings_9 ( // @[PoolingController.scala 23:31]
    .io_pixel1(Max_Poolings_9_io_pixel1),
    .io_pixel2(Max_Poolings_9_io_pixel2),
    .io_pixel3(Max_Poolings_9_io_pixel3),
    .io_pixel4(Max_Poolings_9_io_pixel4),
    .io_f_max(Max_Poolings_9_io_f_max)
  );
  Max_Pooling Max_Poolings_10 ( // @[PoolingController.scala 23:31]
    .io_pixel1(Max_Poolings_10_io_pixel1),
    .io_pixel2(Max_Poolings_10_io_pixel2),
    .io_pixel3(Max_Poolings_10_io_pixel3),
    .io_pixel4(Max_Poolings_10_io_pixel4),
    .io_f_max(Max_Poolings_10_io_f_max)
  );
  Max_Pooling Max_Poolings_11 ( // @[PoolingController.scala 23:31]
    .io_pixel1(Max_Poolings_11_io_pixel1),
    .io_pixel2(Max_Poolings_11_io_pixel2),
    .io_pixel3(Max_Poolings_11_io_pixel3),
    .io_pixel4(Max_Poolings_11_io_pixel4),
    .io_f_max(Max_Poolings_11_io_f_max)
  );
  Max_Pooling Max_Poolings_12 ( // @[PoolingController.scala 23:31]
    .io_pixel1(Max_Poolings_12_io_pixel1),
    .io_pixel2(Max_Poolings_12_io_pixel2),
    .io_pixel3(Max_Poolings_12_io_pixel3),
    .io_pixel4(Max_Poolings_12_io_pixel4),
    .io_f_max(Max_Poolings_12_io_f_max)
  );
  Max_Pooling Max_Poolings_13 ( // @[PoolingController.scala 23:31]
    .io_pixel1(Max_Poolings_13_io_pixel1),
    .io_pixel2(Max_Poolings_13_io_pixel2),
    .io_pixel3(Max_Poolings_13_io_pixel3),
    .io_pixel4(Max_Poolings_13_io_pixel4),
    .io_f_max(Max_Poolings_13_io_f_max)
  );
  Max_Pooling Max_Poolings_14 ( // @[PoolingController.scala 23:31]
    .io_pixel1(Max_Poolings_14_io_pixel1),
    .io_pixel2(Max_Poolings_14_io_pixel2),
    .io_pixel3(Max_Poolings_14_io_pixel3),
    .io_pixel4(Max_Poolings_14_io_pixel4),
    .io_f_max(Max_Poolings_14_io_f_max)
  );
  Max_Pooling Max_Poolings_15 ( // @[PoolingController.scala 23:31]
    .io_pixel1(Max_Poolings_15_io_pixel1),
    .io_pixel2(Max_Poolings_15_io_pixel2),
    .io_pixel3(Max_Poolings_15_io_pixel3),
    .io_pixel4(Max_Poolings_15_io_pixel4),
    .io_f_max(Max_Poolings_15_io_f_max)
  );
  assign io_single_out_0 = Max_Poolings_0_io_f_max; // @[PoolingController.scala 47:23]
  assign io_single_out_1 = Max_Poolings_1_io_f_max; // @[PoolingController.scala 47:23]
  assign io_single_out_2 = Max_Poolings_2_io_f_max; // @[PoolingController.scala 47:23]
  assign io_single_out_3 = Max_Poolings_3_io_f_max; // @[PoolingController.scala 47:23]
  assign io_single_out_4 = Max_Poolings_4_io_f_max; // @[PoolingController.scala 47:23]
  assign io_single_out_5 = Max_Poolings_5_io_f_max; // @[PoolingController.scala 47:23]
  assign io_single_out_6 = Max_Poolings_6_io_f_max; // @[PoolingController.scala 47:23]
  assign io_single_out_7 = Max_Poolings_7_io_f_max; // @[PoolingController.scala 47:23]
  assign io_single_out_8 = Max_Poolings_8_io_f_max; // @[PoolingController.scala 47:23]
  assign io_single_out_9 = Max_Poolings_9_io_f_max; // @[PoolingController.scala 47:23]
  assign io_single_out_10 = Max_Poolings_10_io_f_max; // @[PoolingController.scala 47:23]
  assign io_single_out_11 = Max_Poolings_11_io_f_max; // @[PoolingController.scala 47:23]
  assign io_single_out_12 = Max_Poolings_12_io_f_max; // @[PoolingController.scala 47:23]
  assign io_single_out_13 = Max_Poolings_13_io_f_max; // @[PoolingController.scala 47:23]
  assign io_single_out_14 = Max_Poolings_14_io_f_max; // @[PoolingController.scala 47:23]
  assign io_single_out_15 = Max_Poolings_15_io_f_max; // @[PoolingController.scala 47:23]
  assign Max_Poolings_0_io_pixel1 = values_0; // @[PoolingController.scala 43:33]
  assign Max_Poolings_0_io_pixel2 = values_1; // @[PoolingController.scala 44:33]
  assign Max_Poolings_0_io_pixel3 = values_2; // @[PoolingController.scala 45:33]
  assign Max_Poolings_0_io_pixel4 = values_3; // @[PoolingController.scala 46:33]
  assign Max_Poolings_1_io_pixel1 = values_4; // @[PoolingController.scala 43:33]
  assign Max_Poolings_1_io_pixel2 = values_5; // @[PoolingController.scala 44:33]
  assign Max_Poolings_1_io_pixel3 = values_6; // @[PoolingController.scala 45:33]
  assign Max_Poolings_1_io_pixel4 = values_7; // @[PoolingController.scala 46:33]
  assign Max_Poolings_2_io_pixel1 = values_8; // @[PoolingController.scala 43:33]
  assign Max_Poolings_2_io_pixel2 = values_9; // @[PoolingController.scala 44:33]
  assign Max_Poolings_2_io_pixel3 = values_10; // @[PoolingController.scala 45:33]
  assign Max_Poolings_2_io_pixel4 = values_11; // @[PoolingController.scala 46:33]
  assign Max_Poolings_3_io_pixel1 = values_12; // @[PoolingController.scala 43:33]
  assign Max_Poolings_3_io_pixel2 = values_13; // @[PoolingController.scala 44:33]
  assign Max_Poolings_3_io_pixel3 = values_14; // @[PoolingController.scala 45:33]
  assign Max_Poolings_3_io_pixel4 = values_15; // @[PoolingController.scala 46:33]
  assign Max_Poolings_4_io_pixel1 = values_16; // @[PoolingController.scala 43:33]
  assign Max_Poolings_4_io_pixel2 = values_17; // @[PoolingController.scala 44:33]
  assign Max_Poolings_4_io_pixel3 = values_18; // @[PoolingController.scala 45:33]
  assign Max_Poolings_4_io_pixel4 = values_19; // @[PoolingController.scala 46:33]
  assign Max_Poolings_5_io_pixel1 = values_20; // @[PoolingController.scala 43:33]
  assign Max_Poolings_5_io_pixel2 = values_21; // @[PoolingController.scala 44:33]
  assign Max_Poolings_5_io_pixel3 = values_22; // @[PoolingController.scala 45:33]
  assign Max_Poolings_5_io_pixel4 = values_23; // @[PoolingController.scala 46:33]
  assign Max_Poolings_6_io_pixel1 = values_24; // @[PoolingController.scala 43:33]
  assign Max_Poolings_6_io_pixel2 = values_25; // @[PoolingController.scala 44:33]
  assign Max_Poolings_6_io_pixel3 = values_26; // @[PoolingController.scala 45:33]
  assign Max_Poolings_6_io_pixel4 = values_27; // @[PoolingController.scala 46:33]
  assign Max_Poolings_7_io_pixel1 = values_28; // @[PoolingController.scala 43:33]
  assign Max_Poolings_7_io_pixel2 = values_29; // @[PoolingController.scala 44:33]
  assign Max_Poolings_7_io_pixel3 = values_30; // @[PoolingController.scala 45:33]
  assign Max_Poolings_7_io_pixel4 = values_31; // @[PoolingController.scala 46:33]
  assign Max_Poolings_8_io_pixel1 = values_32; // @[PoolingController.scala 43:33]
  assign Max_Poolings_8_io_pixel2 = values_33; // @[PoolingController.scala 44:33]
  assign Max_Poolings_8_io_pixel3 = values_34; // @[PoolingController.scala 45:33]
  assign Max_Poolings_8_io_pixel4 = values_35; // @[PoolingController.scala 46:33]
  assign Max_Poolings_9_io_pixel1 = values_36; // @[PoolingController.scala 43:33]
  assign Max_Poolings_9_io_pixel2 = values_37; // @[PoolingController.scala 44:33]
  assign Max_Poolings_9_io_pixel3 = values_38; // @[PoolingController.scala 45:33]
  assign Max_Poolings_9_io_pixel4 = values_39; // @[PoolingController.scala 46:33]
  assign Max_Poolings_10_io_pixel1 = values_40; // @[PoolingController.scala 43:33]
  assign Max_Poolings_10_io_pixel2 = values_41; // @[PoolingController.scala 44:33]
  assign Max_Poolings_10_io_pixel3 = values_42; // @[PoolingController.scala 45:33]
  assign Max_Poolings_10_io_pixel4 = values_43; // @[PoolingController.scala 46:33]
  assign Max_Poolings_11_io_pixel1 = values_44; // @[PoolingController.scala 43:33]
  assign Max_Poolings_11_io_pixel2 = values_45; // @[PoolingController.scala 44:33]
  assign Max_Poolings_11_io_pixel3 = values_46; // @[PoolingController.scala 45:33]
  assign Max_Poolings_11_io_pixel4 = values_47; // @[PoolingController.scala 46:33]
  assign Max_Poolings_12_io_pixel1 = values_48; // @[PoolingController.scala 43:33]
  assign Max_Poolings_12_io_pixel2 = values_49; // @[PoolingController.scala 44:33]
  assign Max_Poolings_12_io_pixel3 = values_50; // @[PoolingController.scala 45:33]
  assign Max_Poolings_12_io_pixel4 = values_51; // @[PoolingController.scala 46:33]
  assign Max_Poolings_13_io_pixel1 = values_52; // @[PoolingController.scala 43:33]
  assign Max_Poolings_13_io_pixel2 = values_53; // @[PoolingController.scala 44:33]
  assign Max_Poolings_13_io_pixel3 = values_54; // @[PoolingController.scala 45:33]
  assign Max_Poolings_13_io_pixel4 = values_55; // @[PoolingController.scala 46:33]
  assign Max_Poolings_14_io_pixel1 = values_56; // @[PoolingController.scala 43:33]
  assign Max_Poolings_14_io_pixel2 = values_57; // @[PoolingController.scala 44:33]
  assign Max_Poolings_14_io_pixel3 = values_58; // @[PoolingController.scala 45:33]
  assign Max_Poolings_14_io_pixel4 = values_59; // @[PoolingController.scala 46:33]
  assign Max_Poolings_15_io_pixel1 = values_60; // @[PoolingController.scala 43:33]
  assign Max_Poolings_15_io_pixel2 = values_61; // @[PoolingController.scala 44:33]
  assign Max_Poolings_15_io_pixel3 = values_62; // @[PoolingController.scala 45:33]
  assign Max_Poolings_15_io_pixel4 = values_63; // @[PoolingController.scala 46:33]
  always @(posedge clock) begin
    values_0 <= io_InputMatrix_0; // @[PoolingController.scala 36:29]
    values_1 <= io_InputMatrix_1; // @[PoolingController.scala 36:29]
    values_2 <= io_InputMatrix_8; // @[PoolingController.scala 36:29]
    values_3 <= io_InputMatrix_9; // @[PoolingController.scala 36:29]
    values_4 <= io_InputMatrix_2; // @[PoolingController.scala 36:29]
    values_5 <= io_InputMatrix_3; // @[PoolingController.scala 36:29]
    values_6 <= io_InputMatrix_10; // @[PoolingController.scala 36:29]
    values_7 <= io_InputMatrix_11; // @[PoolingController.scala 36:29]
    values_8 <= io_InputMatrix_4; // @[PoolingController.scala 36:29]
    values_9 <= io_InputMatrix_5; // @[PoolingController.scala 36:29]
    values_10 <= io_InputMatrix_12; // @[PoolingController.scala 36:29]
    values_11 <= io_InputMatrix_13; // @[PoolingController.scala 36:29]
    values_12 <= io_InputMatrix_6; // @[PoolingController.scala 36:29]
    values_13 <= io_InputMatrix_7; // @[PoolingController.scala 36:29]
    values_14 <= io_InputMatrix_14; // @[PoolingController.scala 36:29]
    values_15 <= io_InputMatrix_15; // @[PoolingController.scala 36:29]
    values_16 <= io_InputMatrix_16; // @[PoolingController.scala 36:29]
    values_17 <= io_InputMatrix_17; // @[PoolingController.scala 36:29]
    values_18 <= io_InputMatrix_24; // @[PoolingController.scala 36:29]
    values_19 <= io_InputMatrix_25; // @[PoolingController.scala 36:29]
    values_20 <= io_InputMatrix_18; // @[PoolingController.scala 36:29]
    values_21 <= io_InputMatrix_19; // @[PoolingController.scala 36:29]
    values_22 <= io_InputMatrix_26; // @[PoolingController.scala 36:29]
    values_23 <= io_InputMatrix_27; // @[PoolingController.scala 36:29]
    values_24 <= io_InputMatrix_20; // @[PoolingController.scala 36:29]
    values_25 <= io_InputMatrix_21; // @[PoolingController.scala 36:29]
    values_26 <= io_InputMatrix_28; // @[PoolingController.scala 36:29]
    values_27 <= io_InputMatrix_29; // @[PoolingController.scala 36:29]
    values_28 <= io_InputMatrix_22; // @[PoolingController.scala 36:29]
    values_29 <= io_InputMatrix_23; // @[PoolingController.scala 36:29]
    values_30 <= io_InputMatrix_30; // @[PoolingController.scala 36:29]
    values_31 <= io_InputMatrix_31; // @[PoolingController.scala 36:29]
    values_32 <= io_InputMatrix_32; // @[PoolingController.scala 36:29]
    values_33 <= io_InputMatrix_33; // @[PoolingController.scala 36:29]
    values_34 <= io_InputMatrix_40; // @[PoolingController.scala 36:29]
    values_35 <= io_InputMatrix_41; // @[PoolingController.scala 36:29]
    values_36 <= io_InputMatrix_34; // @[PoolingController.scala 36:29]
    values_37 <= io_InputMatrix_35; // @[PoolingController.scala 36:29]
    values_38 <= io_InputMatrix_42; // @[PoolingController.scala 36:29]
    values_39 <= io_InputMatrix_43; // @[PoolingController.scala 36:29]
    values_40 <= io_InputMatrix_36; // @[PoolingController.scala 36:29]
    values_41 <= io_InputMatrix_37; // @[PoolingController.scala 36:29]
    values_42 <= io_InputMatrix_44; // @[PoolingController.scala 36:29]
    values_43 <= io_InputMatrix_45; // @[PoolingController.scala 36:29]
    values_44 <= io_InputMatrix_38; // @[PoolingController.scala 36:29]
    values_45 <= io_InputMatrix_39; // @[PoolingController.scala 36:29]
    values_46 <= io_InputMatrix_46; // @[PoolingController.scala 36:29]
    values_47 <= io_InputMatrix_47; // @[PoolingController.scala 36:29]
    values_48 <= io_InputMatrix_48; // @[PoolingController.scala 36:29]
    values_49 <= io_InputMatrix_49; // @[PoolingController.scala 36:29]
    values_50 <= io_InputMatrix_56; // @[PoolingController.scala 36:29]
    values_51 <= io_InputMatrix_57; // @[PoolingController.scala 36:29]
    values_52 <= io_InputMatrix_50; // @[PoolingController.scala 36:29]
    values_53 <= io_InputMatrix_51; // @[PoolingController.scala 36:29]
    values_54 <= io_InputMatrix_58; // @[PoolingController.scala 36:29]
    values_55 <= io_InputMatrix_59; // @[PoolingController.scala 36:29]
    values_56 <= io_InputMatrix_52; // @[PoolingController.scala 36:29]
    values_57 <= io_InputMatrix_53; // @[PoolingController.scala 36:29]
    values_58 <= io_InputMatrix_60; // @[PoolingController.scala 36:29]
    values_59 <= io_InputMatrix_61; // @[PoolingController.scala 36:29]
    values_60 <= io_InputMatrix_54; // @[PoolingController.scala 36:29]
    values_61 <= io_InputMatrix_55; // @[PoolingController.scala 36:29]
    values_62 <= io_InputMatrix_62; // @[PoolingController.scala 36:29]
    values_63 <= io_InputMatrix_63; // @[PoolingController.scala 36:29]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  values_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  values_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  values_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  values_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  values_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  values_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  values_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  values_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  values_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  values_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  values_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  values_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  values_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  values_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  values_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  values_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  values_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  values_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  values_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  values_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  values_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  values_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  values_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  values_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  values_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  values_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  values_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  values_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  values_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  values_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  values_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  values_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  values_32 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  values_33 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  values_34 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  values_35 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  values_36 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  values_37 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  values_38 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  values_39 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  values_40 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  values_41 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  values_42 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  values_43 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  values_44 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  values_45 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  values_46 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  values_47 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  values_48 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  values_49 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  values_50 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  values_51 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  values_52 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  values_53 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  values_54 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  values_55 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  values_56 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  values_57 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  values_58 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  values_59 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  values_60 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  values_61 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  values_62 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  values_63 = _RAND_63[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FP_multiply_sum_64(
  input  [31:0] io_in_a_0,
  input  [31:0] io_in_a_1,
  input  [31:0] io_in_a_2,
  input  [31:0] io_in_a_3,
  input  [31:0] io_in_a_4,
  input  [31:0] io_in_a_5,
  input  [31:0] io_in_a_6,
  input  [31:0] io_in_a_7,
  input  [31:0] io_in_a_8,
  input  [31:0] io_in_a_9,
  input  [31:0] io_in_a_10,
  input  [31:0] io_in_a_11,
  input  [31:0] io_in_a_12,
  input  [31:0] io_in_a_13,
  input  [31:0] io_in_a_14,
  input  [31:0] io_in_a_15,
  input  [31:0] io_in_b_0,
  input  [31:0] io_in_b_1,
  input  [31:0] io_in_b_2,
  input  [31:0] io_in_b_3,
  input  [31:0] io_in_b_4,
  input  [31:0] io_in_b_5,
  input  [31:0] io_in_b_6,
  input  [31:0] io_in_b_7,
  input  [31:0] io_in_b_8,
  input  [31:0] io_in_b_9,
  input  [31:0] io_in_b_10,
  input  [31:0] io_in_b_11,
  input  [31:0] io_in_b_12,
  input  [31:0] io_in_b_13,
  input  [31:0] io_in_b_14,
  input  [31:0] io_in_b_15,
  output [31:0] io_out_s
);
  wire [31:0] FP_multipliers_0_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_0_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_0_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_1_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_1_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_1_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_2_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_2_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_2_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_3_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_3_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_3_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_4_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_4_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_4_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_5_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_5_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_5_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_6_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_6_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_6_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_7_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_7_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_7_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_8_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_8_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_8_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_9_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_9_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_9_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_10_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_10_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_10_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_11_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_11_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_11_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_12_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_12_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_12_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_13_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_13_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_13_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_14_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_14_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_14_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_15_io_in_a; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_15_io_in_b; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_multipliers_15_io_out_s; // @[FPArithmetic.scala 623:33]
  wire [31:0] FP_adders_0_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_0_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_0_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_1_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_1_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_1_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_2_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_2_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_2_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_3_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_3_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_3_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_4_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_4_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_4_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_5_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_5_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_5_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_6_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_6_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_6_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_7_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_7_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_7_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_8_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_8_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_8_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_9_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_9_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_9_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_10_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_10_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_10_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_11_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_11_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_11_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_12_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_12_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_12_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_13_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_13_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_13_io_out_s; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_14_io_in_a; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_14_io_in_b; // @[FPArithmetic.scala 630:28]
  wire [31:0] FP_adders_14_io_out_s; // @[FPArithmetic.scala 630:28]
  FP_multiplier FP_multipliers_0 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_0_io_in_a),
    .io_in_b(FP_multipliers_0_io_in_b),
    .io_out_s(FP_multipliers_0_io_out_s)
  );
  FP_multiplier FP_multipliers_1 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_1_io_in_a),
    .io_in_b(FP_multipliers_1_io_in_b),
    .io_out_s(FP_multipliers_1_io_out_s)
  );
  FP_multiplier FP_multipliers_2 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_2_io_in_a),
    .io_in_b(FP_multipliers_2_io_in_b),
    .io_out_s(FP_multipliers_2_io_out_s)
  );
  FP_multiplier FP_multipliers_3 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_3_io_in_a),
    .io_in_b(FP_multipliers_3_io_in_b),
    .io_out_s(FP_multipliers_3_io_out_s)
  );
  FP_multiplier FP_multipliers_4 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_4_io_in_a),
    .io_in_b(FP_multipliers_4_io_in_b),
    .io_out_s(FP_multipliers_4_io_out_s)
  );
  FP_multiplier FP_multipliers_5 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_5_io_in_a),
    .io_in_b(FP_multipliers_5_io_in_b),
    .io_out_s(FP_multipliers_5_io_out_s)
  );
  FP_multiplier FP_multipliers_6 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_6_io_in_a),
    .io_in_b(FP_multipliers_6_io_in_b),
    .io_out_s(FP_multipliers_6_io_out_s)
  );
  FP_multiplier FP_multipliers_7 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_7_io_in_a),
    .io_in_b(FP_multipliers_7_io_in_b),
    .io_out_s(FP_multipliers_7_io_out_s)
  );
  FP_multiplier FP_multipliers_8 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_8_io_in_a),
    .io_in_b(FP_multipliers_8_io_in_b),
    .io_out_s(FP_multipliers_8_io_out_s)
  );
  FP_multiplier FP_multipliers_9 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_9_io_in_a),
    .io_in_b(FP_multipliers_9_io_in_b),
    .io_out_s(FP_multipliers_9_io_out_s)
  );
  FP_multiplier FP_multipliers_10 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_10_io_in_a),
    .io_in_b(FP_multipliers_10_io_in_b),
    .io_out_s(FP_multipliers_10_io_out_s)
  );
  FP_multiplier FP_multipliers_11 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_11_io_in_a),
    .io_in_b(FP_multipliers_11_io_in_b),
    .io_out_s(FP_multipliers_11_io_out_s)
  );
  FP_multiplier FP_multipliers_12 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_12_io_in_a),
    .io_in_b(FP_multipliers_12_io_in_b),
    .io_out_s(FP_multipliers_12_io_out_s)
  );
  FP_multiplier FP_multipliers_13 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_13_io_in_a),
    .io_in_b(FP_multipliers_13_io_in_b),
    .io_out_s(FP_multipliers_13_io_out_s)
  );
  FP_multiplier FP_multipliers_14 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_14_io_in_a),
    .io_in_b(FP_multipliers_14_io_in_b),
    .io_out_s(FP_multipliers_14_io_out_s)
  );
  FP_multiplier FP_multipliers_15 ( // @[FPArithmetic.scala 623:33]
    .io_in_a(FP_multipliers_15_io_in_a),
    .io_in_b(FP_multipliers_15_io_in_b),
    .io_out_s(FP_multipliers_15_io_out_s)
  );
  FP_adder FP_adders_0 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_0_io_in_a),
    .io_in_b(FP_adders_0_io_in_b),
    .io_out_s(FP_adders_0_io_out_s)
  );
  FP_adder FP_adders_1 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_1_io_in_a),
    .io_in_b(FP_adders_1_io_in_b),
    .io_out_s(FP_adders_1_io_out_s)
  );
  FP_adder FP_adders_2 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_2_io_in_a),
    .io_in_b(FP_adders_2_io_in_b),
    .io_out_s(FP_adders_2_io_out_s)
  );
  FP_adder FP_adders_3 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_3_io_in_a),
    .io_in_b(FP_adders_3_io_in_b),
    .io_out_s(FP_adders_3_io_out_s)
  );
  FP_adder FP_adders_4 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_4_io_in_a),
    .io_in_b(FP_adders_4_io_in_b),
    .io_out_s(FP_adders_4_io_out_s)
  );
  FP_adder FP_adders_5 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_5_io_in_a),
    .io_in_b(FP_adders_5_io_in_b),
    .io_out_s(FP_adders_5_io_out_s)
  );
  FP_adder FP_adders_6 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_6_io_in_a),
    .io_in_b(FP_adders_6_io_in_b),
    .io_out_s(FP_adders_6_io_out_s)
  );
  FP_adder FP_adders_7 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_7_io_in_a),
    .io_in_b(FP_adders_7_io_in_b),
    .io_out_s(FP_adders_7_io_out_s)
  );
  FP_adder FP_adders_8 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_8_io_in_a),
    .io_in_b(FP_adders_8_io_in_b),
    .io_out_s(FP_adders_8_io_out_s)
  );
  FP_adder FP_adders_9 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_9_io_in_a),
    .io_in_b(FP_adders_9_io_in_b),
    .io_out_s(FP_adders_9_io_out_s)
  );
  FP_adder FP_adders_10 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_10_io_in_a),
    .io_in_b(FP_adders_10_io_in_b),
    .io_out_s(FP_adders_10_io_out_s)
  );
  FP_adder FP_adders_11 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_11_io_in_a),
    .io_in_b(FP_adders_11_io_in_b),
    .io_out_s(FP_adders_11_io_out_s)
  );
  FP_adder FP_adders_12 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_12_io_in_a),
    .io_in_b(FP_adders_12_io_in_b),
    .io_out_s(FP_adders_12_io_out_s)
  );
  FP_adder FP_adders_13 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_13_io_in_a),
    .io_in_b(FP_adders_13_io_in_b),
    .io_out_s(FP_adders_13_io_out_s)
  );
  FP_adder FP_adders_14 ( // @[FPArithmetic.scala 630:28]
    .io_in_a(FP_adders_14_io_in_a),
    .io_in_b(FP_adders_14_io_in_b),
    .io_out_s(FP_adders_14_io_out_s)
  );
  assign io_out_s = FP_adders_14_io_out_s; // @[FPArithmetic.scala 693:14]
  assign FP_multipliers_0_io_in_a = io_in_a_0; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_0_io_in_b = io_in_b_0; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_1_io_in_a = io_in_a_1; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_1_io_in_b = io_in_b_1; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_2_io_in_a = io_in_a_2; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_2_io_in_b = io_in_b_2; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_3_io_in_a = io_in_a_3; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_3_io_in_b = io_in_b_3; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_4_io_in_a = io_in_a_4; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_4_io_in_b = io_in_b_4; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_5_io_in_a = io_in_a_5; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_5_io_in_b = io_in_b_5; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_6_io_in_a = io_in_a_6; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_6_io_in_b = io_in_b_6; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_7_io_in_a = io_in_a_7; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_7_io_in_b = io_in_b_7; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_8_io_in_a = io_in_a_8; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_8_io_in_b = io_in_b_8; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_9_io_in_a = io_in_a_9; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_9_io_in_b = io_in_b_9; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_10_io_in_a = io_in_a_10; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_10_io_in_b = io_in_b_10; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_11_io_in_a = io_in_a_11; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_11_io_in_b = io_in_b_11; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_12_io_in_a = io_in_a_12; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_12_io_in_b = io_in_b_12; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_13_io_in_a = io_in_a_13; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_13_io_in_b = io_in_b_13; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_14_io_in_a = io_in_a_14; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_14_io_in_b = io_in_b_14; // @[FPArithmetic.scala 637:33]
  assign FP_multipliers_15_io_in_a = io_in_a_15; // @[FPArithmetic.scala 636:33]
  assign FP_multipliers_15_io_in_b = io_in_b_15; // @[FPArithmetic.scala 637:33]
  assign FP_adders_0_io_in_a = FP_multipliers_0_io_out_s; // @[FPArithmetic.scala 655:41]
  assign FP_adders_0_io_in_b = FP_multipliers_1_io_out_s; // @[FPArithmetic.scala 656:41]
  assign FP_adders_1_io_in_a = FP_multipliers_2_io_out_s; // @[FPArithmetic.scala 655:41]
  assign FP_adders_1_io_in_b = FP_multipliers_3_io_out_s; // @[FPArithmetic.scala 656:41]
  assign FP_adders_2_io_in_a = FP_multipliers_4_io_out_s; // @[FPArithmetic.scala 655:41]
  assign FP_adders_2_io_in_b = FP_multipliers_5_io_out_s; // @[FPArithmetic.scala 656:41]
  assign FP_adders_3_io_in_a = FP_multipliers_6_io_out_s; // @[FPArithmetic.scala 655:41]
  assign FP_adders_3_io_in_b = FP_multipliers_7_io_out_s; // @[FPArithmetic.scala 656:41]
  assign FP_adders_4_io_in_a = FP_multipliers_8_io_out_s; // @[FPArithmetic.scala 655:41]
  assign FP_adders_4_io_in_b = FP_multipliers_9_io_out_s; // @[FPArithmetic.scala 656:41]
  assign FP_adders_5_io_in_a = FP_multipliers_10_io_out_s; // @[FPArithmetic.scala 655:41]
  assign FP_adders_5_io_in_b = FP_multipliers_11_io_out_s; // @[FPArithmetic.scala 656:41]
  assign FP_adders_6_io_in_a = FP_multipliers_12_io_out_s; // @[FPArithmetic.scala 655:41]
  assign FP_adders_6_io_in_b = FP_multipliers_13_io_out_s; // @[FPArithmetic.scala 656:41]
  assign FP_adders_7_io_in_a = FP_multipliers_14_io_out_s; // @[FPArithmetic.scala 655:41]
  assign FP_adders_7_io_in_b = FP_multipliers_15_io_out_s; // @[FPArithmetic.scala 656:41]
  assign FP_adders_8_io_in_a = FP_adders_0_io_out_s; // @[FPArithmetic.scala 681:43]
  assign FP_adders_8_io_in_b = FP_adders_1_io_out_s; // @[FPArithmetic.scala 682:43]
  assign FP_adders_9_io_in_a = FP_adders_2_io_out_s; // @[FPArithmetic.scala 681:43]
  assign FP_adders_9_io_in_b = FP_adders_3_io_out_s; // @[FPArithmetic.scala 682:43]
  assign FP_adders_10_io_in_a = FP_adders_4_io_out_s; // @[FPArithmetic.scala 681:43]
  assign FP_adders_10_io_in_b = FP_adders_5_io_out_s; // @[FPArithmetic.scala 682:43]
  assign FP_adders_11_io_in_a = FP_adders_6_io_out_s; // @[FPArithmetic.scala 681:43]
  assign FP_adders_11_io_in_b = FP_adders_7_io_out_s; // @[FPArithmetic.scala 682:43]
  assign FP_adders_12_io_in_a = FP_adders_8_io_out_s; // @[FPArithmetic.scala 681:43]
  assign FP_adders_12_io_in_b = FP_adders_9_io_out_s; // @[FPArithmetic.scala 682:43]
  assign FP_adders_13_io_in_a = FP_adders_10_io_out_s; // @[FPArithmetic.scala 681:43]
  assign FP_adders_13_io_in_b = FP_adders_11_io_out_s; // @[FPArithmetic.scala 682:43]
  assign FP_adders_14_io_in_a = FP_adders_12_io_out_s; // @[FPArithmetic.scala 681:43]
  assign FP_adders_14_io_in_b = FP_adders_13_io_out_s; // @[FPArithmetic.scala 682:43]
endmodule
module FC(
  input  [31:0] io_matB_0,
  input  [31:0] io_matB_1,
  input  [31:0] io_matB_2,
  input  [31:0] io_matB_3,
  input  [31:0] io_matB_4,
  input  [31:0] io_matB_5,
  input  [31:0] io_matB_6,
  input  [31:0] io_matB_7,
  input  [31:0] io_matB_8,
  input  [31:0] io_matB_9,
  input  [31:0] io_matB_10,
  input  [31:0] io_matB_11,
  input  [31:0] io_matB_12,
  input  [31:0] io_matB_13,
  input  [31:0] io_matB_14,
  input  [31:0] io_matB_15,
  output [31:0] io_fC_out_0,
  output [31:0] io_fC_out_1,
  output [31:0] io_fC_out_2,
  output [31:0] io_fC_out_3,
  output [31:0] io_fC_out_4,
  output [31:0] io_fC_out_5,
  output [31:0] io_fC_out_6,
  output [31:0] io_fC_out_7,
  output [31:0] io_fC_out_8,
  output [31:0] io_fC_out_9
);
  wire [31:0] mul_io_in_a_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_a_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_a_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_a_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_a_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_a_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_a_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_a_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_a_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_a_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_a_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_a_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_a_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_a_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_a_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_a_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_b_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_b_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_b_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_b_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_b_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_b_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_b_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_b_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_b_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_b_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_b_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_b_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_b_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_b_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_b_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_in_b_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_io_out_s; // @[FCLayer.scala 18:23]
  wire [31:0] fp_adder_io_in_a; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_io_in_b; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_io_out_s; // @[FCLayer.scala 23:28]
  wire [31:0] mul_1_io_in_a_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_a_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_a_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_a_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_a_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_a_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_a_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_a_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_a_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_a_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_a_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_a_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_a_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_a_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_a_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_a_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_b_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_b_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_b_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_b_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_b_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_b_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_b_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_b_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_b_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_b_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_b_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_b_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_b_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_b_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_b_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_in_b_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_1_io_out_s; // @[FCLayer.scala 18:23]
  wire [31:0] fp_adder_1_io_in_a; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_1_io_in_b; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_1_io_out_s; // @[FCLayer.scala 23:28]
  wire [31:0] mul_2_io_in_a_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_a_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_a_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_a_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_a_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_a_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_a_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_a_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_a_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_a_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_a_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_a_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_a_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_a_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_a_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_a_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_b_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_b_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_b_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_b_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_b_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_b_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_b_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_b_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_b_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_b_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_b_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_b_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_b_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_b_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_b_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_in_b_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_2_io_out_s; // @[FCLayer.scala 18:23]
  wire [31:0] fp_adder_2_io_in_a; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_2_io_in_b; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_2_io_out_s; // @[FCLayer.scala 23:28]
  wire [31:0] mul_3_io_in_a_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_a_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_a_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_a_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_a_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_a_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_a_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_a_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_a_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_a_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_a_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_a_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_a_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_a_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_a_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_a_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_b_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_b_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_b_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_b_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_b_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_b_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_b_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_b_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_b_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_b_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_b_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_b_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_b_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_b_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_b_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_in_b_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_3_io_out_s; // @[FCLayer.scala 18:23]
  wire [31:0] fp_adder_3_io_in_a; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_3_io_in_b; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_3_io_out_s; // @[FCLayer.scala 23:28]
  wire [31:0] mul_4_io_in_a_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_a_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_a_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_a_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_a_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_a_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_a_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_a_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_a_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_a_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_a_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_a_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_a_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_a_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_a_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_a_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_b_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_b_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_b_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_b_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_b_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_b_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_b_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_b_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_b_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_b_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_b_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_b_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_b_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_b_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_b_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_in_b_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_4_io_out_s; // @[FCLayer.scala 18:23]
  wire [31:0] fp_adder_4_io_in_a; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_4_io_in_b; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_4_io_out_s; // @[FCLayer.scala 23:28]
  wire [31:0] mul_5_io_in_a_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_a_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_a_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_a_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_a_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_a_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_a_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_a_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_a_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_a_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_a_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_a_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_a_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_a_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_a_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_a_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_b_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_b_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_b_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_b_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_b_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_b_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_b_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_b_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_b_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_b_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_b_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_b_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_b_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_b_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_b_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_in_b_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_5_io_out_s; // @[FCLayer.scala 18:23]
  wire [31:0] fp_adder_5_io_in_a; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_5_io_in_b; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_5_io_out_s; // @[FCLayer.scala 23:28]
  wire [31:0] mul_6_io_in_a_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_a_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_a_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_a_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_a_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_a_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_a_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_a_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_a_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_a_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_a_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_a_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_a_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_a_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_a_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_a_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_b_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_b_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_b_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_b_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_b_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_b_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_b_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_b_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_b_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_b_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_b_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_b_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_b_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_b_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_b_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_in_b_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_6_io_out_s; // @[FCLayer.scala 18:23]
  wire [31:0] fp_adder_6_io_in_a; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_6_io_in_b; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_6_io_out_s; // @[FCLayer.scala 23:28]
  wire [31:0] mul_7_io_in_a_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_a_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_a_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_a_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_a_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_a_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_a_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_a_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_a_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_a_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_a_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_a_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_a_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_a_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_a_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_a_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_b_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_b_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_b_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_b_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_b_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_b_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_b_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_b_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_b_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_b_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_b_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_b_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_b_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_b_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_b_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_in_b_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_7_io_out_s; // @[FCLayer.scala 18:23]
  wire [31:0] fp_adder_7_io_in_a; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_7_io_in_b; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_7_io_out_s; // @[FCLayer.scala 23:28]
  wire [31:0] mul_8_io_in_a_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_a_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_a_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_a_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_a_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_a_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_a_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_a_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_a_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_a_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_a_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_a_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_a_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_a_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_a_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_a_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_b_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_b_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_b_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_b_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_b_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_b_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_b_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_b_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_b_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_b_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_b_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_b_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_b_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_b_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_b_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_in_b_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_8_io_out_s; // @[FCLayer.scala 18:23]
  wire [31:0] fp_adder_8_io_in_a; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_8_io_in_b; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_8_io_out_s; // @[FCLayer.scala 23:28]
  wire [31:0] mul_9_io_in_a_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_a_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_a_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_a_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_a_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_a_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_a_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_a_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_a_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_a_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_a_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_a_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_a_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_a_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_a_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_a_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_b_0; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_b_1; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_b_2; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_b_3; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_b_4; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_b_5; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_b_6; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_b_7; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_b_8; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_b_9; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_b_10; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_b_11; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_b_12; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_b_13; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_b_14; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_in_b_15; // @[FCLayer.scala 18:23]
  wire [31:0] mul_9_io_out_s; // @[FCLayer.scala 18:23]
  wire [31:0] fp_adder_9_io_in_a; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_9_io_in_b; // @[FCLayer.scala 23:28]
  wire [31:0] fp_adder_9_io_out_s; // @[FCLayer.scala 23:28]
  FP_multiply_sum_64 mul ( // @[FCLayer.scala 18:23]
    .io_in_a_0(mul_io_in_a_0),
    .io_in_a_1(mul_io_in_a_1),
    .io_in_a_2(mul_io_in_a_2),
    .io_in_a_3(mul_io_in_a_3),
    .io_in_a_4(mul_io_in_a_4),
    .io_in_a_5(mul_io_in_a_5),
    .io_in_a_6(mul_io_in_a_6),
    .io_in_a_7(mul_io_in_a_7),
    .io_in_a_8(mul_io_in_a_8),
    .io_in_a_9(mul_io_in_a_9),
    .io_in_a_10(mul_io_in_a_10),
    .io_in_a_11(mul_io_in_a_11),
    .io_in_a_12(mul_io_in_a_12),
    .io_in_a_13(mul_io_in_a_13),
    .io_in_a_14(mul_io_in_a_14),
    .io_in_a_15(mul_io_in_a_15),
    .io_in_b_0(mul_io_in_b_0),
    .io_in_b_1(mul_io_in_b_1),
    .io_in_b_2(mul_io_in_b_2),
    .io_in_b_3(mul_io_in_b_3),
    .io_in_b_4(mul_io_in_b_4),
    .io_in_b_5(mul_io_in_b_5),
    .io_in_b_6(mul_io_in_b_6),
    .io_in_b_7(mul_io_in_b_7),
    .io_in_b_8(mul_io_in_b_8),
    .io_in_b_9(mul_io_in_b_9),
    .io_in_b_10(mul_io_in_b_10),
    .io_in_b_11(mul_io_in_b_11),
    .io_in_b_12(mul_io_in_b_12),
    .io_in_b_13(mul_io_in_b_13),
    .io_in_b_14(mul_io_in_b_14),
    .io_in_b_15(mul_io_in_b_15),
    .io_out_s(mul_io_out_s)
  );
  FP_adder fp_adder ( // @[FCLayer.scala 23:28]
    .io_in_a(fp_adder_io_in_a),
    .io_in_b(fp_adder_io_in_b),
    .io_out_s(fp_adder_io_out_s)
  );
  FP_multiply_sum_64 mul_1 ( // @[FCLayer.scala 18:23]
    .io_in_a_0(mul_1_io_in_a_0),
    .io_in_a_1(mul_1_io_in_a_1),
    .io_in_a_2(mul_1_io_in_a_2),
    .io_in_a_3(mul_1_io_in_a_3),
    .io_in_a_4(mul_1_io_in_a_4),
    .io_in_a_5(mul_1_io_in_a_5),
    .io_in_a_6(mul_1_io_in_a_6),
    .io_in_a_7(mul_1_io_in_a_7),
    .io_in_a_8(mul_1_io_in_a_8),
    .io_in_a_9(mul_1_io_in_a_9),
    .io_in_a_10(mul_1_io_in_a_10),
    .io_in_a_11(mul_1_io_in_a_11),
    .io_in_a_12(mul_1_io_in_a_12),
    .io_in_a_13(mul_1_io_in_a_13),
    .io_in_a_14(mul_1_io_in_a_14),
    .io_in_a_15(mul_1_io_in_a_15),
    .io_in_b_0(mul_1_io_in_b_0),
    .io_in_b_1(mul_1_io_in_b_1),
    .io_in_b_2(mul_1_io_in_b_2),
    .io_in_b_3(mul_1_io_in_b_3),
    .io_in_b_4(mul_1_io_in_b_4),
    .io_in_b_5(mul_1_io_in_b_5),
    .io_in_b_6(mul_1_io_in_b_6),
    .io_in_b_7(mul_1_io_in_b_7),
    .io_in_b_8(mul_1_io_in_b_8),
    .io_in_b_9(mul_1_io_in_b_9),
    .io_in_b_10(mul_1_io_in_b_10),
    .io_in_b_11(mul_1_io_in_b_11),
    .io_in_b_12(mul_1_io_in_b_12),
    .io_in_b_13(mul_1_io_in_b_13),
    .io_in_b_14(mul_1_io_in_b_14),
    .io_in_b_15(mul_1_io_in_b_15),
    .io_out_s(mul_1_io_out_s)
  );
  FP_adder fp_adder_1 ( // @[FCLayer.scala 23:28]
    .io_in_a(fp_adder_1_io_in_a),
    .io_in_b(fp_adder_1_io_in_b),
    .io_out_s(fp_adder_1_io_out_s)
  );
  FP_multiply_sum_64 mul_2 ( // @[FCLayer.scala 18:23]
    .io_in_a_0(mul_2_io_in_a_0),
    .io_in_a_1(mul_2_io_in_a_1),
    .io_in_a_2(mul_2_io_in_a_2),
    .io_in_a_3(mul_2_io_in_a_3),
    .io_in_a_4(mul_2_io_in_a_4),
    .io_in_a_5(mul_2_io_in_a_5),
    .io_in_a_6(mul_2_io_in_a_6),
    .io_in_a_7(mul_2_io_in_a_7),
    .io_in_a_8(mul_2_io_in_a_8),
    .io_in_a_9(mul_2_io_in_a_9),
    .io_in_a_10(mul_2_io_in_a_10),
    .io_in_a_11(mul_2_io_in_a_11),
    .io_in_a_12(mul_2_io_in_a_12),
    .io_in_a_13(mul_2_io_in_a_13),
    .io_in_a_14(mul_2_io_in_a_14),
    .io_in_a_15(mul_2_io_in_a_15),
    .io_in_b_0(mul_2_io_in_b_0),
    .io_in_b_1(mul_2_io_in_b_1),
    .io_in_b_2(mul_2_io_in_b_2),
    .io_in_b_3(mul_2_io_in_b_3),
    .io_in_b_4(mul_2_io_in_b_4),
    .io_in_b_5(mul_2_io_in_b_5),
    .io_in_b_6(mul_2_io_in_b_6),
    .io_in_b_7(mul_2_io_in_b_7),
    .io_in_b_8(mul_2_io_in_b_8),
    .io_in_b_9(mul_2_io_in_b_9),
    .io_in_b_10(mul_2_io_in_b_10),
    .io_in_b_11(mul_2_io_in_b_11),
    .io_in_b_12(mul_2_io_in_b_12),
    .io_in_b_13(mul_2_io_in_b_13),
    .io_in_b_14(mul_2_io_in_b_14),
    .io_in_b_15(mul_2_io_in_b_15),
    .io_out_s(mul_2_io_out_s)
  );
  FP_adder fp_adder_2 ( // @[FCLayer.scala 23:28]
    .io_in_a(fp_adder_2_io_in_a),
    .io_in_b(fp_adder_2_io_in_b),
    .io_out_s(fp_adder_2_io_out_s)
  );
  FP_multiply_sum_64 mul_3 ( // @[FCLayer.scala 18:23]
    .io_in_a_0(mul_3_io_in_a_0),
    .io_in_a_1(mul_3_io_in_a_1),
    .io_in_a_2(mul_3_io_in_a_2),
    .io_in_a_3(mul_3_io_in_a_3),
    .io_in_a_4(mul_3_io_in_a_4),
    .io_in_a_5(mul_3_io_in_a_5),
    .io_in_a_6(mul_3_io_in_a_6),
    .io_in_a_7(mul_3_io_in_a_7),
    .io_in_a_8(mul_3_io_in_a_8),
    .io_in_a_9(mul_3_io_in_a_9),
    .io_in_a_10(mul_3_io_in_a_10),
    .io_in_a_11(mul_3_io_in_a_11),
    .io_in_a_12(mul_3_io_in_a_12),
    .io_in_a_13(mul_3_io_in_a_13),
    .io_in_a_14(mul_3_io_in_a_14),
    .io_in_a_15(mul_3_io_in_a_15),
    .io_in_b_0(mul_3_io_in_b_0),
    .io_in_b_1(mul_3_io_in_b_1),
    .io_in_b_2(mul_3_io_in_b_2),
    .io_in_b_3(mul_3_io_in_b_3),
    .io_in_b_4(mul_3_io_in_b_4),
    .io_in_b_5(mul_3_io_in_b_5),
    .io_in_b_6(mul_3_io_in_b_6),
    .io_in_b_7(mul_3_io_in_b_7),
    .io_in_b_8(mul_3_io_in_b_8),
    .io_in_b_9(mul_3_io_in_b_9),
    .io_in_b_10(mul_3_io_in_b_10),
    .io_in_b_11(mul_3_io_in_b_11),
    .io_in_b_12(mul_3_io_in_b_12),
    .io_in_b_13(mul_3_io_in_b_13),
    .io_in_b_14(mul_3_io_in_b_14),
    .io_in_b_15(mul_3_io_in_b_15),
    .io_out_s(mul_3_io_out_s)
  );
  FP_adder fp_adder_3 ( // @[FCLayer.scala 23:28]
    .io_in_a(fp_adder_3_io_in_a),
    .io_in_b(fp_adder_3_io_in_b),
    .io_out_s(fp_adder_3_io_out_s)
  );
  FP_multiply_sum_64 mul_4 ( // @[FCLayer.scala 18:23]
    .io_in_a_0(mul_4_io_in_a_0),
    .io_in_a_1(mul_4_io_in_a_1),
    .io_in_a_2(mul_4_io_in_a_2),
    .io_in_a_3(mul_4_io_in_a_3),
    .io_in_a_4(mul_4_io_in_a_4),
    .io_in_a_5(mul_4_io_in_a_5),
    .io_in_a_6(mul_4_io_in_a_6),
    .io_in_a_7(mul_4_io_in_a_7),
    .io_in_a_8(mul_4_io_in_a_8),
    .io_in_a_9(mul_4_io_in_a_9),
    .io_in_a_10(mul_4_io_in_a_10),
    .io_in_a_11(mul_4_io_in_a_11),
    .io_in_a_12(mul_4_io_in_a_12),
    .io_in_a_13(mul_4_io_in_a_13),
    .io_in_a_14(mul_4_io_in_a_14),
    .io_in_a_15(mul_4_io_in_a_15),
    .io_in_b_0(mul_4_io_in_b_0),
    .io_in_b_1(mul_4_io_in_b_1),
    .io_in_b_2(mul_4_io_in_b_2),
    .io_in_b_3(mul_4_io_in_b_3),
    .io_in_b_4(mul_4_io_in_b_4),
    .io_in_b_5(mul_4_io_in_b_5),
    .io_in_b_6(mul_4_io_in_b_6),
    .io_in_b_7(mul_4_io_in_b_7),
    .io_in_b_8(mul_4_io_in_b_8),
    .io_in_b_9(mul_4_io_in_b_9),
    .io_in_b_10(mul_4_io_in_b_10),
    .io_in_b_11(mul_4_io_in_b_11),
    .io_in_b_12(mul_4_io_in_b_12),
    .io_in_b_13(mul_4_io_in_b_13),
    .io_in_b_14(mul_4_io_in_b_14),
    .io_in_b_15(mul_4_io_in_b_15),
    .io_out_s(mul_4_io_out_s)
  );
  FP_adder fp_adder_4 ( // @[FCLayer.scala 23:28]
    .io_in_a(fp_adder_4_io_in_a),
    .io_in_b(fp_adder_4_io_in_b),
    .io_out_s(fp_adder_4_io_out_s)
  );
  FP_multiply_sum_64 mul_5 ( // @[FCLayer.scala 18:23]
    .io_in_a_0(mul_5_io_in_a_0),
    .io_in_a_1(mul_5_io_in_a_1),
    .io_in_a_2(mul_5_io_in_a_2),
    .io_in_a_3(mul_5_io_in_a_3),
    .io_in_a_4(mul_5_io_in_a_4),
    .io_in_a_5(mul_5_io_in_a_5),
    .io_in_a_6(mul_5_io_in_a_6),
    .io_in_a_7(mul_5_io_in_a_7),
    .io_in_a_8(mul_5_io_in_a_8),
    .io_in_a_9(mul_5_io_in_a_9),
    .io_in_a_10(mul_5_io_in_a_10),
    .io_in_a_11(mul_5_io_in_a_11),
    .io_in_a_12(mul_5_io_in_a_12),
    .io_in_a_13(mul_5_io_in_a_13),
    .io_in_a_14(mul_5_io_in_a_14),
    .io_in_a_15(mul_5_io_in_a_15),
    .io_in_b_0(mul_5_io_in_b_0),
    .io_in_b_1(mul_5_io_in_b_1),
    .io_in_b_2(mul_5_io_in_b_2),
    .io_in_b_3(mul_5_io_in_b_3),
    .io_in_b_4(mul_5_io_in_b_4),
    .io_in_b_5(mul_5_io_in_b_5),
    .io_in_b_6(mul_5_io_in_b_6),
    .io_in_b_7(mul_5_io_in_b_7),
    .io_in_b_8(mul_5_io_in_b_8),
    .io_in_b_9(mul_5_io_in_b_9),
    .io_in_b_10(mul_5_io_in_b_10),
    .io_in_b_11(mul_5_io_in_b_11),
    .io_in_b_12(mul_5_io_in_b_12),
    .io_in_b_13(mul_5_io_in_b_13),
    .io_in_b_14(mul_5_io_in_b_14),
    .io_in_b_15(mul_5_io_in_b_15),
    .io_out_s(mul_5_io_out_s)
  );
  FP_adder fp_adder_5 ( // @[FCLayer.scala 23:28]
    .io_in_a(fp_adder_5_io_in_a),
    .io_in_b(fp_adder_5_io_in_b),
    .io_out_s(fp_adder_5_io_out_s)
  );
  FP_multiply_sum_64 mul_6 ( // @[FCLayer.scala 18:23]
    .io_in_a_0(mul_6_io_in_a_0),
    .io_in_a_1(mul_6_io_in_a_1),
    .io_in_a_2(mul_6_io_in_a_2),
    .io_in_a_3(mul_6_io_in_a_3),
    .io_in_a_4(mul_6_io_in_a_4),
    .io_in_a_5(mul_6_io_in_a_5),
    .io_in_a_6(mul_6_io_in_a_6),
    .io_in_a_7(mul_6_io_in_a_7),
    .io_in_a_8(mul_6_io_in_a_8),
    .io_in_a_9(mul_6_io_in_a_9),
    .io_in_a_10(mul_6_io_in_a_10),
    .io_in_a_11(mul_6_io_in_a_11),
    .io_in_a_12(mul_6_io_in_a_12),
    .io_in_a_13(mul_6_io_in_a_13),
    .io_in_a_14(mul_6_io_in_a_14),
    .io_in_a_15(mul_6_io_in_a_15),
    .io_in_b_0(mul_6_io_in_b_0),
    .io_in_b_1(mul_6_io_in_b_1),
    .io_in_b_2(mul_6_io_in_b_2),
    .io_in_b_3(mul_6_io_in_b_3),
    .io_in_b_4(mul_6_io_in_b_4),
    .io_in_b_5(mul_6_io_in_b_5),
    .io_in_b_6(mul_6_io_in_b_6),
    .io_in_b_7(mul_6_io_in_b_7),
    .io_in_b_8(mul_6_io_in_b_8),
    .io_in_b_9(mul_6_io_in_b_9),
    .io_in_b_10(mul_6_io_in_b_10),
    .io_in_b_11(mul_6_io_in_b_11),
    .io_in_b_12(mul_6_io_in_b_12),
    .io_in_b_13(mul_6_io_in_b_13),
    .io_in_b_14(mul_6_io_in_b_14),
    .io_in_b_15(mul_6_io_in_b_15),
    .io_out_s(mul_6_io_out_s)
  );
  FP_adder fp_adder_6 ( // @[FCLayer.scala 23:28]
    .io_in_a(fp_adder_6_io_in_a),
    .io_in_b(fp_adder_6_io_in_b),
    .io_out_s(fp_adder_6_io_out_s)
  );
  FP_multiply_sum_64 mul_7 ( // @[FCLayer.scala 18:23]
    .io_in_a_0(mul_7_io_in_a_0),
    .io_in_a_1(mul_7_io_in_a_1),
    .io_in_a_2(mul_7_io_in_a_2),
    .io_in_a_3(mul_7_io_in_a_3),
    .io_in_a_4(mul_7_io_in_a_4),
    .io_in_a_5(mul_7_io_in_a_5),
    .io_in_a_6(mul_7_io_in_a_6),
    .io_in_a_7(mul_7_io_in_a_7),
    .io_in_a_8(mul_7_io_in_a_8),
    .io_in_a_9(mul_7_io_in_a_9),
    .io_in_a_10(mul_7_io_in_a_10),
    .io_in_a_11(mul_7_io_in_a_11),
    .io_in_a_12(mul_7_io_in_a_12),
    .io_in_a_13(mul_7_io_in_a_13),
    .io_in_a_14(mul_7_io_in_a_14),
    .io_in_a_15(mul_7_io_in_a_15),
    .io_in_b_0(mul_7_io_in_b_0),
    .io_in_b_1(mul_7_io_in_b_1),
    .io_in_b_2(mul_7_io_in_b_2),
    .io_in_b_3(mul_7_io_in_b_3),
    .io_in_b_4(mul_7_io_in_b_4),
    .io_in_b_5(mul_7_io_in_b_5),
    .io_in_b_6(mul_7_io_in_b_6),
    .io_in_b_7(mul_7_io_in_b_7),
    .io_in_b_8(mul_7_io_in_b_8),
    .io_in_b_9(mul_7_io_in_b_9),
    .io_in_b_10(mul_7_io_in_b_10),
    .io_in_b_11(mul_7_io_in_b_11),
    .io_in_b_12(mul_7_io_in_b_12),
    .io_in_b_13(mul_7_io_in_b_13),
    .io_in_b_14(mul_7_io_in_b_14),
    .io_in_b_15(mul_7_io_in_b_15),
    .io_out_s(mul_7_io_out_s)
  );
  FP_adder fp_adder_7 ( // @[FCLayer.scala 23:28]
    .io_in_a(fp_adder_7_io_in_a),
    .io_in_b(fp_adder_7_io_in_b),
    .io_out_s(fp_adder_7_io_out_s)
  );
  FP_multiply_sum_64 mul_8 ( // @[FCLayer.scala 18:23]
    .io_in_a_0(mul_8_io_in_a_0),
    .io_in_a_1(mul_8_io_in_a_1),
    .io_in_a_2(mul_8_io_in_a_2),
    .io_in_a_3(mul_8_io_in_a_3),
    .io_in_a_4(mul_8_io_in_a_4),
    .io_in_a_5(mul_8_io_in_a_5),
    .io_in_a_6(mul_8_io_in_a_6),
    .io_in_a_7(mul_8_io_in_a_7),
    .io_in_a_8(mul_8_io_in_a_8),
    .io_in_a_9(mul_8_io_in_a_9),
    .io_in_a_10(mul_8_io_in_a_10),
    .io_in_a_11(mul_8_io_in_a_11),
    .io_in_a_12(mul_8_io_in_a_12),
    .io_in_a_13(mul_8_io_in_a_13),
    .io_in_a_14(mul_8_io_in_a_14),
    .io_in_a_15(mul_8_io_in_a_15),
    .io_in_b_0(mul_8_io_in_b_0),
    .io_in_b_1(mul_8_io_in_b_1),
    .io_in_b_2(mul_8_io_in_b_2),
    .io_in_b_3(mul_8_io_in_b_3),
    .io_in_b_4(mul_8_io_in_b_4),
    .io_in_b_5(mul_8_io_in_b_5),
    .io_in_b_6(mul_8_io_in_b_6),
    .io_in_b_7(mul_8_io_in_b_7),
    .io_in_b_8(mul_8_io_in_b_8),
    .io_in_b_9(mul_8_io_in_b_9),
    .io_in_b_10(mul_8_io_in_b_10),
    .io_in_b_11(mul_8_io_in_b_11),
    .io_in_b_12(mul_8_io_in_b_12),
    .io_in_b_13(mul_8_io_in_b_13),
    .io_in_b_14(mul_8_io_in_b_14),
    .io_in_b_15(mul_8_io_in_b_15),
    .io_out_s(mul_8_io_out_s)
  );
  FP_adder fp_adder_8 ( // @[FCLayer.scala 23:28]
    .io_in_a(fp_adder_8_io_in_a),
    .io_in_b(fp_adder_8_io_in_b),
    .io_out_s(fp_adder_8_io_out_s)
  );
  FP_multiply_sum_64 mul_9 ( // @[FCLayer.scala 18:23]
    .io_in_a_0(mul_9_io_in_a_0),
    .io_in_a_1(mul_9_io_in_a_1),
    .io_in_a_2(mul_9_io_in_a_2),
    .io_in_a_3(mul_9_io_in_a_3),
    .io_in_a_4(mul_9_io_in_a_4),
    .io_in_a_5(mul_9_io_in_a_5),
    .io_in_a_6(mul_9_io_in_a_6),
    .io_in_a_7(mul_9_io_in_a_7),
    .io_in_a_8(mul_9_io_in_a_8),
    .io_in_a_9(mul_9_io_in_a_9),
    .io_in_a_10(mul_9_io_in_a_10),
    .io_in_a_11(mul_9_io_in_a_11),
    .io_in_a_12(mul_9_io_in_a_12),
    .io_in_a_13(mul_9_io_in_a_13),
    .io_in_a_14(mul_9_io_in_a_14),
    .io_in_a_15(mul_9_io_in_a_15),
    .io_in_b_0(mul_9_io_in_b_0),
    .io_in_b_1(mul_9_io_in_b_1),
    .io_in_b_2(mul_9_io_in_b_2),
    .io_in_b_3(mul_9_io_in_b_3),
    .io_in_b_4(mul_9_io_in_b_4),
    .io_in_b_5(mul_9_io_in_b_5),
    .io_in_b_6(mul_9_io_in_b_6),
    .io_in_b_7(mul_9_io_in_b_7),
    .io_in_b_8(mul_9_io_in_b_8),
    .io_in_b_9(mul_9_io_in_b_9),
    .io_in_b_10(mul_9_io_in_b_10),
    .io_in_b_11(mul_9_io_in_b_11),
    .io_in_b_12(mul_9_io_in_b_12),
    .io_in_b_13(mul_9_io_in_b_13),
    .io_in_b_14(mul_9_io_in_b_14),
    .io_in_b_15(mul_9_io_in_b_15),
    .io_out_s(mul_9_io_out_s)
  );
  FP_adder fp_adder_9 ( // @[FCLayer.scala 23:28]
    .io_in_a(fp_adder_9_io_in_a),
    .io_in_b(fp_adder_9_io_in_b),
    .io_out_s(fp_adder_9_io_out_s)
  );
  assign io_fC_out_0 = fp_adder_io_out_s; // @[FCLayer.scala 26:20]
  assign io_fC_out_1 = fp_adder_1_io_out_s; // @[FCLayer.scala 26:20]
  assign io_fC_out_2 = fp_adder_2_io_out_s; // @[FCLayer.scala 26:20]
  assign io_fC_out_3 = fp_adder_3_io_out_s; // @[FCLayer.scala 26:20]
  assign io_fC_out_4 = fp_adder_4_io_out_s; // @[FCLayer.scala 26:20]
  assign io_fC_out_5 = fp_adder_5_io_out_s; // @[FCLayer.scala 26:20]
  assign io_fC_out_6 = fp_adder_6_io_out_s; // @[FCLayer.scala 26:20]
  assign io_fC_out_7 = fp_adder_7_io_out_s; // @[FCLayer.scala 26:20]
  assign io_fC_out_8 = fp_adder_8_io_out_s; // @[FCLayer.scala 26:20]
  assign io_fC_out_9 = fp_adder_9_io_out_s; // @[FCLayer.scala 26:20]
  assign mul_io_in_a_0 = 32'h3dccccc0; // @[FCLayer.scala 20:24]
  assign mul_io_in_a_1 = 32'h3dccccc0; // @[FCLayer.scala 20:24]
  assign mul_io_in_a_2 = 32'h3e6147a8; // @[FCLayer.scala 20:24]
  assign mul_io_in_a_3 = 32'h3dccccc0; // @[FCLayer.scala 20:24]
  assign mul_io_in_a_4 = 32'h3de147a0; // @[FCLayer.scala 20:24]
  assign mul_io_in_a_5 = 32'h3de147a0; // @[FCLayer.scala 20:24]
  assign mul_io_in_a_6 = 32'h3de147a0; // @[FCLayer.scala 20:24]
  assign mul_io_in_a_7 = 32'h3f8020c4; // @[FCLayer.scala 20:24]
  assign mul_io_in_a_8 = 32'h3e4cccc8; // @[FCLayer.scala 20:24]
  assign mul_io_in_a_9 = 32'h3f333332; // @[FCLayer.scala 20:24]
  assign mul_io_in_a_10 = 32'h3d8f5c20; // @[FCLayer.scala 20:24]
  assign mul_io_in_a_11 = 32'h3dccccc0; // @[FCLayer.scala 20:24]
  assign mul_io_in_a_12 = 32'h3e6b8518; // @[FCLayer.scala 20:24]
  assign mul_io_in_a_13 = 32'h3e75c288; // @[FCLayer.scala 20:24]
  assign mul_io_in_a_14 = 32'h3e6b8518; // @[FCLayer.scala 20:24]
  assign mul_io_in_a_15 = 32'h3e6147a8; // @[FCLayer.scala 20:24]
  assign mul_io_in_b_0 = io_matB_0; // @[FCLayer.scala 21:24]
  assign mul_io_in_b_1 = io_matB_1; // @[FCLayer.scala 21:24]
  assign mul_io_in_b_2 = io_matB_2; // @[FCLayer.scala 21:24]
  assign mul_io_in_b_3 = io_matB_3; // @[FCLayer.scala 21:24]
  assign mul_io_in_b_4 = io_matB_4; // @[FCLayer.scala 21:24]
  assign mul_io_in_b_5 = io_matB_5; // @[FCLayer.scala 21:24]
  assign mul_io_in_b_6 = io_matB_6; // @[FCLayer.scala 21:24]
  assign mul_io_in_b_7 = io_matB_7; // @[FCLayer.scala 21:24]
  assign mul_io_in_b_8 = io_matB_8; // @[FCLayer.scala 21:24]
  assign mul_io_in_b_9 = io_matB_9; // @[FCLayer.scala 21:24]
  assign mul_io_in_b_10 = io_matB_10; // @[FCLayer.scala 21:24]
  assign mul_io_in_b_11 = io_matB_11; // @[FCLayer.scala 21:24]
  assign mul_io_in_b_12 = io_matB_12; // @[FCLayer.scala 21:24]
  assign mul_io_in_b_13 = io_matB_13; // @[FCLayer.scala 21:24]
  assign mul_io_in_b_14 = io_matB_14; // @[FCLayer.scala 21:24]
  assign mul_io_in_b_15 = io_matB_15; // @[FCLayer.scala 21:24]
  assign fp_adder_io_in_a = mul_io_out_s; // @[FCLayer.scala 24:24]
  assign fp_adder_io_in_b = 32'h3f800000; // @[FCLayer.scala 25:24]
  assign mul_1_io_in_a_0 = 32'h3df5c280; // @[FCLayer.scala 20:24]
  assign mul_1_io_in_a_1 = 32'h3e75c288; // @[FCLayer.scala 20:24]
  assign mul_1_io_in_a_2 = 32'h3de147a0; // @[FCLayer.scala 20:24]
  assign mul_1_io_in_a_3 = 32'h3f63d70a; // @[FCLayer.scala 20:24]
  assign mul_1_io_in_a_4 = 32'h40333333; // @[FCLayer.scala 20:24]
  assign mul_1_io_in_a_5 = 32'h3e6147a8; // @[FCLayer.scala 20:24]
  assign mul_1_io_in_a_6 = 32'h40933333; // @[FCLayer.scala 20:24]
  assign mul_1_io_in_a_7 = 32'h3f8a3d70; // @[FCLayer.scala 20:24]
  assign mul_1_io_in_a_8 = 32'h3eae1478; // @[FCLayer.scala 20:24]
  assign mul_1_io_in_a_9 = 32'h4007ae14; // @[FCLayer.scala 20:24]
  assign mul_1_io_in_a_10 = 32'h3f23d70a; // @[FCLayer.scala 20:24]
  assign mul_1_io_in_a_11 = 32'h3d23d700; // @[FCLayer.scala 20:24]
  assign mul_1_io_in_a_12 = 32'h3eae1478; // @[FCLayer.scala 20:24]
  assign mul_1_io_in_a_13 = 32'h3f9d70a3; // @[FCLayer.scala 20:24]
  assign mul_1_io_in_a_14 = 32'h40066666; // @[FCLayer.scala 20:24]
  assign mul_1_io_in_a_15 = 32'h3f8ccccc; // @[FCLayer.scala 20:24]
  assign mul_1_io_in_b_0 = io_matB_0; // @[FCLayer.scala 21:24]
  assign mul_1_io_in_b_1 = io_matB_1; // @[FCLayer.scala 21:24]
  assign mul_1_io_in_b_2 = io_matB_2; // @[FCLayer.scala 21:24]
  assign mul_1_io_in_b_3 = io_matB_3; // @[FCLayer.scala 21:24]
  assign mul_1_io_in_b_4 = io_matB_4; // @[FCLayer.scala 21:24]
  assign mul_1_io_in_b_5 = io_matB_5; // @[FCLayer.scala 21:24]
  assign mul_1_io_in_b_6 = io_matB_6; // @[FCLayer.scala 21:24]
  assign mul_1_io_in_b_7 = io_matB_7; // @[FCLayer.scala 21:24]
  assign mul_1_io_in_b_8 = io_matB_8; // @[FCLayer.scala 21:24]
  assign mul_1_io_in_b_9 = io_matB_9; // @[FCLayer.scala 21:24]
  assign mul_1_io_in_b_10 = io_matB_10; // @[FCLayer.scala 21:24]
  assign mul_1_io_in_b_11 = io_matB_11; // @[FCLayer.scala 21:24]
  assign mul_1_io_in_b_12 = io_matB_12; // @[FCLayer.scala 21:24]
  assign mul_1_io_in_b_13 = io_matB_13; // @[FCLayer.scala 21:24]
  assign mul_1_io_in_b_14 = io_matB_14; // @[FCLayer.scala 21:24]
  assign mul_1_io_in_b_15 = io_matB_15; // @[FCLayer.scala 21:24]
  assign fp_adder_1_io_in_a = mul_1_io_out_s; // @[FCLayer.scala 24:24]
  assign fp_adder_1_io_in_b = 32'h3e4cccc8; // @[FCLayer.scala 25:24]
  assign mul_2_io_in_a_0 = 32'h3f9c28f5; // @[FCLayer.scala 20:24]
  assign mul_2_io_in_a_1 = 32'h40466666; // @[FCLayer.scala 20:24]
  assign mul_2_io_in_a_2 = 32'h40c3851e; // @[FCLayer.scala 20:24]
  assign mul_2_io_in_a_3 = 32'h4111c28f; // @[FCLayer.scala 20:24]
  assign mul_2_io_in_a_4 = 32'h40070a3d; // @[FCLayer.scala 20:24]
  assign mul_2_io_in_a_5 = 32'h3f8020c4; // @[FCLayer.scala 20:24]
  assign mul_2_io_in_a_6 = 32'h404ccccc; // @[FCLayer.scala 20:24]
  assign mul_2_io_in_a_7 = 32'h40d66666; // @[FCLayer.scala 20:24]
  assign mul_2_io_in_a_8 = 32'h41011eb8; // @[FCLayer.scala 20:24]
  assign mul_2_io_in_a_9 = 32'h40066666; // @[FCLayer.scala 20:24]
  assign mul_2_io_in_a_10 = 32'h3f9d70a3; // @[FCLayer.scala 20:24]
  assign mul_2_io_in_a_11 = 32'h404f5c28; // @[FCLayer.scala 20:24]
  assign mul_2_io_in_a_12 = 32'h3f9d70a3; // @[FCLayer.scala 20:24]
  assign mul_2_io_in_a_13 = 32'h404e147a; // @[FCLayer.scala 20:24]
  assign mul_2_io_in_a_14 = 32'h40a3d70a; // @[FCLayer.scala 20:24]
  assign mul_2_io_in_a_15 = 32'h404f5c28; // @[FCLayer.scala 20:24]
  assign mul_2_io_in_b_0 = io_matB_0; // @[FCLayer.scala 21:24]
  assign mul_2_io_in_b_1 = io_matB_1; // @[FCLayer.scala 21:24]
  assign mul_2_io_in_b_2 = io_matB_2; // @[FCLayer.scala 21:24]
  assign mul_2_io_in_b_3 = io_matB_3; // @[FCLayer.scala 21:24]
  assign mul_2_io_in_b_4 = io_matB_4; // @[FCLayer.scala 21:24]
  assign mul_2_io_in_b_5 = io_matB_5; // @[FCLayer.scala 21:24]
  assign mul_2_io_in_b_6 = io_matB_6; // @[FCLayer.scala 21:24]
  assign mul_2_io_in_b_7 = io_matB_7; // @[FCLayer.scala 21:24]
  assign mul_2_io_in_b_8 = io_matB_8; // @[FCLayer.scala 21:24]
  assign mul_2_io_in_b_9 = io_matB_9; // @[FCLayer.scala 21:24]
  assign mul_2_io_in_b_10 = io_matB_10; // @[FCLayer.scala 21:24]
  assign mul_2_io_in_b_11 = io_matB_11; // @[FCLayer.scala 21:24]
  assign mul_2_io_in_b_12 = io_matB_12; // @[FCLayer.scala 21:24]
  assign mul_2_io_in_b_13 = io_matB_13; // @[FCLayer.scala 21:24]
  assign mul_2_io_in_b_14 = io_matB_14; // @[FCLayer.scala 21:24]
  assign mul_2_io_in_b_15 = io_matB_15; // @[FCLayer.scala 21:24]
  assign fp_adder_2_io_in_a = mul_2_io_out_s; // @[FCLayer.scala 24:24]
  assign fp_adder_2_io_in_b = 32'h3dccccc0; // @[FCLayer.scala 25:24]
  assign mul_3_io_in_a_0 = 32'h3f8e147a; // @[FCLayer.scala 20:24]
  assign mul_3_io_in_a_1 = 32'h3f63d70a; // @[FCLayer.scala 20:24]
  assign mul_3_io_in_a_2 = 32'h40333333; // @[FCLayer.scala 20:24]
  assign mul_3_io_in_a_3 = 32'h400e147a; // @[FCLayer.scala 20:24]
  assign mul_3_io_in_a_4 = 32'h40933333; // @[FCLayer.scala 20:24]
  assign mul_3_io_in_a_5 = 32'h3f8a3d70; // @[FCLayer.scala 20:24]
  assign mul_3_io_in_a_6 = 32'h4015c28f; // @[FCLayer.scala 20:24]
  assign mul_3_io_in_a_7 = 32'h4007ae14; // @[FCLayer.scala 20:24]
  assign mul_3_io_in_a_8 = 32'h40f47ae1; // @[FCLayer.scala 20:24]
  assign mul_3_io_in_a_9 = 32'h4110a3d7; // @[FCLayer.scala 20:24]
  assign mul_3_io_in_a_10 = 32'h4015c28f; // @[FCLayer.scala 20:24]
  assign mul_3_io_in_a_11 = 32'h3f9d70a3; // @[FCLayer.scala 20:24]
  assign mul_3_io_in_a_12 = 32'h40066666; // @[FCLayer.scala 20:24]
  assign mul_3_io_in_a_13 = 32'h3f8ccccc; // @[FCLayer.scala 20:24]
  assign mul_3_io_in_a_14 = 32'h3f9c28f5; // @[FCLayer.scala 20:24]
  assign mul_3_io_in_a_15 = 32'h40466666; // @[FCLayer.scala 20:24]
  assign mul_3_io_in_b_0 = io_matB_0; // @[FCLayer.scala 21:24]
  assign mul_3_io_in_b_1 = io_matB_1; // @[FCLayer.scala 21:24]
  assign mul_3_io_in_b_2 = io_matB_2; // @[FCLayer.scala 21:24]
  assign mul_3_io_in_b_3 = io_matB_3; // @[FCLayer.scala 21:24]
  assign mul_3_io_in_b_4 = io_matB_4; // @[FCLayer.scala 21:24]
  assign mul_3_io_in_b_5 = io_matB_5; // @[FCLayer.scala 21:24]
  assign mul_3_io_in_b_6 = io_matB_6; // @[FCLayer.scala 21:24]
  assign mul_3_io_in_b_7 = io_matB_7; // @[FCLayer.scala 21:24]
  assign mul_3_io_in_b_8 = io_matB_8; // @[FCLayer.scala 21:24]
  assign mul_3_io_in_b_9 = io_matB_9; // @[FCLayer.scala 21:24]
  assign mul_3_io_in_b_10 = io_matB_10; // @[FCLayer.scala 21:24]
  assign mul_3_io_in_b_11 = io_matB_11; // @[FCLayer.scala 21:24]
  assign mul_3_io_in_b_12 = io_matB_12; // @[FCLayer.scala 21:24]
  assign mul_3_io_in_b_13 = io_matB_13; // @[FCLayer.scala 21:24]
  assign mul_3_io_in_b_14 = io_matB_14; // @[FCLayer.scala 21:24]
  assign mul_3_io_in_b_15 = io_matB_15; // @[FCLayer.scala 21:24]
  assign fp_adder_3_io_in_a = mul_3_io_out_s; // @[FCLayer.scala 24:24]
  assign fp_adder_3_io_in_b = 32'h3e999998; // @[FCLayer.scala 25:24]
  assign mul_4_io_in_a_0 = 32'h40c3851e; // @[FCLayer.scala 20:24]
  assign mul_4_io_in_a_1 = 32'h4111c28f; // @[FCLayer.scala 20:24]
  assign mul_4_io_in_a_2 = 32'h40070a3d; // @[FCLayer.scala 20:24]
  assign mul_4_io_in_a_3 = 32'h3f8020c4; // @[FCLayer.scala 20:24]
  assign mul_4_io_in_a_4 = 32'h404ccccc; // @[FCLayer.scala 20:24]
  assign mul_4_io_in_a_5 = 32'h40d66666; // @[FCLayer.scala 20:24]
  assign mul_4_io_in_a_6 = 32'h41011eb8; // @[FCLayer.scala 20:24]
  assign mul_4_io_in_a_7 = 32'h40066666; // @[FCLayer.scala 20:24]
  assign mul_4_io_in_a_8 = 32'h3f9d70a3; // @[FCLayer.scala 20:24]
  assign mul_4_io_in_a_9 = 32'h404f5c28; // @[FCLayer.scala 20:24]
  assign mul_4_io_in_a_10 = 32'h3f9d70a3; // @[FCLayer.scala 20:24]
  assign mul_4_io_in_a_11 = 32'h404e147a; // @[FCLayer.scala 20:24]
  assign mul_4_io_in_a_12 = 32'h40a3d70a; // @[FCLayer.scala 20:24]
  assign mul_4_io_in_a_13 = 32'h404f5c28; // @[FCLayer.scala 20:24]
  assign mul_4_io_in_a_14 = 32'h3f8e147a; // @[FCLayer.scala 20:24]
  assign mul_4_io_in_a_15 = 32'h3f63d70a; // @[FCLayer.scala 20:24]
  assign mul_4_io_in_b_0 = io_matB_0; // @[FCLayer.scala 21:24]
  assign mul_4_io_in_b_1 = io_matB_1; // @[FCLayer.scala 21:24]
  assign mul_4_io_in_b_2 = io_matB_2; // @[FCLayer.scala 21:24]
  assign mul_4_io_in_b_3 = io_matB_3; // @[FCLayer.scala 21:24]
  assign mul_4_io_in_b_4 = io_matB_4; // @[FCLayer.scala 21:24]
  assign mul_4_io_in_b_5 = io_matB_5; // @[FCLayer.scala 21:24]
  assign mul_4_io_in_b_6 = io_matB_6; // @[FCLayer.scala 21:24]
  assign mul_4_io_in_b_7 = io_matB_7; // @[FCLayer.scala 21:24]
  assign mul_4_io_in_b_8 = io_matB_8; // @[FCLayer.scala 21:24]
  assign mul_4_io_in_b_9 = io_matB_9; // @[FCLayer.scala 21:24]
  assign mul_4_io_in_b_10 = io_matB_10; // @[FCLayer.scala 21:24]
  assign mul_4_io_in_b_11 = io_matB_11; // @[FCLayer.scala 21:24]
  assign mul_4_io_in_b_12 = io_matB_12; // @[FCLayer.scala 21:24]
  assign mul_4_io_in_b_13 = io_matB_13; // @[FCLayer.scala 21:24]
  assign mul_4_io_in_b_14 = io_matB_14; // @[FCLayer.scala 21:24]
  assign mul_4_io_in_b_15 = io_matB_15; // @[FCLayer.scala 21:24]
  assign fp_adder_4_io_in_a = mul_4_io_out_s; // @[FCLayer.scala 24:24]
  assign fp_adder_4_io_in_b = 32'h40a00000; // @[FCLayer.scala 25:24]
  assign mul_5_io_in_a_0 = 32'h40333333; // @[FCLayer.scala 20:24]
  assign mul_5_io_in_a_1 = 32'h400e147a; // @[FCLayer.scala 20:24]
  assign mul_5_io_in_a_2 = 32'h40933333; // @[FCLayer.scala 20:24]
  assign mul_5_io_in_a_3 = 32'h3f8a3d70; // @[FCLayer.scala 20:24]
  assign mul_5_io_in_a_4 = 32'h4015c28f; // @[FCLayer.scala 20:24]
  assign mul_5_io_in_a_5 = 32'h4007ae14; // @[FCLayer.scala 20:24]
  assign mul_5_io_in_a_6 = 32'h40f47ae1; // @[FCLayer.scala 20:24]
  assign mul_5_io_in_a_7 = 32'h4110a3d7; // @[FCLayer.scala 20:24]
  assign mul_5_io_in_a_8 = 32'h4015c28f; // @[FCLayer.scala 20:24]
  assign mul_5_io_in_a_9 = 32'h3f9d70a3; // @[FCLayer.scala 20:24]
  assign mul_5_io_in_a_10 = 32'h40066666; // @[FCLayer.scala 20:24]
  assign mul_5_io_in_a_11 = 32'h3f8ccccc; // @[FCLayer.scala 20:24]
  assign mul_5_io_in_a_12 = 32'h3f9c28f5; // @[FCLayer.scala 20:24]
  assign mul_5_io_in_a_13 = 32'h40466666; // @[FCLayer.scala 20:24]
  assign mul_5_io_in_a_14 = 32'h40c3851e; // @[FCLayer.scala 20:24]
  assign mul_5_io_in_a_15 = 32'h4111c28f; // @[FCLayer.scala 20:24]
  assign mul_5_io_in_b_0 = io_matB_0; // @[FCLayer.scala 21:24]
  assign mul_5_io_in_b_1 = io_matB_1; // @[FCLayer.scala 21:24]
  assign mul_5_io_in_b_2 = io_matB_2; // @[FCLayer.scala 21:24]
  assign mul_5_io_in_b_3 = io_matB_3; // @[FCLayer.scala 21:24]
  assign mul_5_io_in_b_4 = io_matB_4; // @[FCLayer.scala 21:24]
  assign mul_5_io_in_b_5 = io_matB_5; // @[FCLayer.scala 21:24]
  assign mul_5_io_in_b_6 = io_matB_6; // @[FCLayer.scala 21:24]
  assign mul_5_io_in_b_7 = io_matB_7; // @[FCLayer.scala 21:24]
  assign mul_5_io_in_b_8 = io_matB_8; // @[FCLayer.scala 21:24]
  assign mul_5_io_in_b_9 = io_matB_9; // @[FCLayer.scala 21:24]
  assign mul_5_io_in_b_10 = io_matB_10; // @[FCLayer.scala 21:24]
  assign mul_5_io_in_b_11 = io_matB_11; // @[FCLayer.scala 21:24]
  assign mul_5_io_in_b_12 = io_matB_12; // @[FCLayer.scala 21:24]
  assign mul_5_io_in_b_13 = io_matB_13; // @[FCLayer.scala 21:24]
  assign mul_5_io_in_b_14 = io_matB_14; // @[FCLayer.scala 21:24]
  assign mul_5_io_in_b_15 = io_matB_15; // @[FCLayer.scala 21:24]
  assign fp_adder_5_io_in_a = mul_5_io_out_s; // @[FCLayer.scala 24:24]
  assign fp_adder_5_io_in_b = 32'h40c00000; // @[FCLayer.scala 25:24]
  assign mul_6_io_in_a_0 = 32'h40070a3d; // @[FCLayer.scala 20:24]
  assign mul_6_io_in_a_1 = 32'h3f8020c4; // @[FCLayer.scala 20:24]
  assign mul_6_io_in_a_2 = 32'h404ccccc; // @[FCLayer.scala 20:24]
  assign mul_6_io_in_a_3 = 32'h40d66666; // @[FCLayer.scala 20:24]
  assign mul_6_io_in_a_4 = 32'h41011eb8; // @[FCLayer.scala 20:24]
  assign mul_6_io_in_a_5 = 32'h40066666; // @[FCLayer.scala 20:24]
  assign mul_6_io_in_a_6 = 32'h3f9d70a3; // @[FCLayer.scala 20:24]
  assign mul_6_io_in_a_7 = 32'h404f5c28; // @[FCLayer.scala 20:24]
  assign mul_6_io_in_a_8 = 32'h3f9d70a3; // @[FCLayer.scala 20:24]
  assign mul_6_io_in_a_9 = 32'h404e147a; // @[FCLayer.scala 20:24]
  assign mul_6_io_in_a_10 = 32'h40a3d70a; // @[FCLayer.scala 20:24]
  assign mul_6_io_in_a_11 = 32'h404f5c28; // @[FCLayer.scala 20:24]
  assign mul_6_io_in_a_12 = 32'h3f8e147a; // @[FCLayer.scala 20:24]
  assign mul_6_io_in_a_13 = 32'h3f63d70a; // @[FCLayer.scala 20:24]
  assign mul_6_io_in_a_14 = 32'h40333333; // @[FCLayer.scala 20:24]
  assign mul_6_io_in_a_15 = 32'h400e147a; // @[FCLayer.scala 20:24]
  assign mul_6_io_in_b_0 = io_matB_0; // @[FCLayer.scala 21:24]
  assign mul_6_io_in_b_1 = io_matB_1; // @[FCLayer.scala 21:24]
  assign mul_6_io_in_b_2 = io_matB_2; // @[FCLayer.scala 21:24]
  assign mul_6_io_in_b_3 = io_matB_3; // @[FCLayer.scala 21:24]
  assign mul_6_io_in_b_4 = io_matB_4; // @[FCLayer.scala 21:24]
  assign mul_6_io_in_b_5 = io_matB_5; // @[FCLayer.scala 21:24]
  assign mul_6_io_in_b_6 = io_matB_6; // @[FCLayer.scala 21:24]
  assign mul_6_io_in_b_7 = io_matB_7; // @[FCLayer.scala 21:24]
  assign mul_6_io_in_b_8 = io_matB_8; // @[FCLayer.scala 21:24]
  assign mul_6_io_in_b_9 = io_matB_9; // @[FCLayer.scala 21:24]
  assign mul_6_io_in_b_10 = io_matB_10; // @[FCLayer.scala 21:24]
  assign mul_6_io_in_b_11 = io_matB_11; // @[FCLayer.scala 21:24]
  assign mul_6_io_in_b_12 = io_matB_12; // @[FCLayer.scala 21:24]
  assign mul_6_io_in_b_13 = io_matB_13; // @[FCLayer.scala 21:24]
  assign mul_6_io_in_b_14 = io_matB_14; // @[FCLayer.scala 21:24]
  assign mul_6_io_in_b_15 = io_matB_15; // @[FCLayer.scala 21:24]
  assign fp_adder_6_io_in_a = mul_6_io_out_s; // @[FCLayer.scala 24:24]
  assign fp_adder_6_io_in_b = 32'h40e00000; // @[FCLayer.scala 25:24]
  assign mul_7_io_in_a_0 = 32'h40933333; // @[FCLayer.scala 20:24]
  assign mul_7_io_in_a_1 = 32'h3f8a3d70; // @[FCLayer.scala 20:24]
  assign mul_7_io_in_a_2 = 32'h4015c28f; // @[FCLayer.scala 20:24]
  assign mul_7_io_in_a_3 = 32'h4007ae14; // @[FCLayer.scala 20:24]
  assign mul_7_io_in_a_4 = 32'h40f47ae1; // @[FCLayer.scala 20:24]
  assign mul_7_io_in_a_5 = 32'h4110a3d7; // @[FCLayer.scala 20:24]
  assign mul_7_io_in_a_6 = 32'h4015c28f; // @[FCLayer.scala 20:24]
  assign mul_7_io_in_a_7 = 32'h3f9d70a3; // @[FCLayer.scala 20:24]
  assign mul_7_io_in_a_8 = 32'h40066666; // @[FCLayer.scala 20:24]
  assign mul_7_io_in_a_9 = 32'h3f8ccccc; // @[FCLayer.scala 20:24]
  assign mul_7_io_in_a_10 = 32'h3f9c28f5; // @[FCLayer.scala 20:24]
  assign mul_7_io_in_a_11 = 32'h40466666; // @[FCLayer.scala 20:24]
  assign mul_7_io_in_a_12 = 32'h40c3851e; // @[FCLayer.scala 20:24]
  assign mul_7_io_in_a_13 = 32'h4111c28f; // @[FCLayer.scala 20:24]
  assign mul_7_io_in_a_14 = 32'h40070a3d; // @[FCLayer.scala 20:24]
  assign mul_7_io_in_a_15 = 32'h3f8020c4; // @[FCLayer.scala 20:24]
  assign mul_7_io_in_b_0 = io_matB_0; // @[FCLayer.scala 21:24]
  assign mul_7_io_in_b_1 = io_matB_1; // @[FCLayer.scala 21:24]
  assign mul_7_io_in_b_2 = io_matB_2; // @[FCLayer.scala 21:24]
  assign mul_7_io_in_b_3 = io_matB_3; // @[FCLayer.scala 21:24]
  assign mul_7_io_in_b_4 = io_matB_4; // @[FCLayer.scala 21:24]
  assign mul_7_io_in_b_5 = io_matB_5; // @[FCLayer.scala 21:24]
  assign mul_7_io_in_b_6 = io_matB_6; // @[FCLayer.scala 21:24]
  assign mul_7_io_in_b_7 = io_matB_7; // @[FCLayer.scala 21:24]
  assign mul_7_io_in_b_8 = io_matB_8; // @[FCLayer.scala 21:24]
  assign mul_7_io_in_b_9 = io_matB_9; // @[FCLayer.scala 21:24]
  assign mul_7_io_in_b_10 = io_matB_10; // @[FCLayer.scala 21:24]
  assign mul_7_io_in_b_11 = io_matB_11; // @[FCLayer.scala 21:24]
  assign mul_7_io_in_b_12 = io_matB_12; // @[FCLayer.scala 21:24]
  assign mul_7_io_in_b_13 = io_matB_13; // @[FCLayer.scala 21:24]
  assign mul_7_io_in_b_14 = io_matB_14; // @[FCLayer.scala 21:24]
  assign mul_7_io_in_b_15 = io_matB_15; // @[FCLayer.scala 21:24]
  assign fp_adder_7_io_in_a = mul_7_io_out_s; // @[FCLayer.scala 24:24]
  assign fp_adder_7_io_in_b = 32'h41000000; // @[FCLayer.scala 25:24]
  assign mul_8_io_in_a_0 = 32'h404ccccc; // @[FCLayer.scala 20:24]
  assign mul_8_io_in_a_1 = 32'h40d66666; // @[FCLayer.scala 20:24]
  assign mul_8_io_in_a_2 = 32'h41011eb8; // @[FCLayer.scala 20:24]
  assign mul_8_io_in_a_3 = 32'h40066666; // @[FCLayer.scala 20:24]
  assign mul_8_io_in_a_4 = 32'h3f9d70a3; // @[FCLayer.scala 20:24]
  assign mul_8_io_in_a_5 = 32'h404f5c28; // @[FCLayer.scala 20:24]
  assign mul_8_io_in_a_6 = 32'h3f9d70a3; // @[FCLayer.scala 20:24]
  assign mul_8_io_in_a_7 = 32'h404e147a; // @[FCLayer.scala 20:24]
  assign mul_8_io_in_a_8 = 32'h40a3d70a; // @[FCLayer.scala 20:24]
  assign mul_8_io_in_a_9 = 32'h404f5c28; // @[FCLayer.scala 20:24]
  assign mul_8_io_in_a_10 = 32'h3f8e147a; // @[FCLayer.scala 20:24]
  assign mul_8_io_in_a_11 = 32'h3f63d70a; // @[FCLayer.scala 20:24]
  assign mul_8_io_in_a_12 = 32'h40333333; // @[FCLayer.scala 20:24]
  assign mul_8_io_in_a_13 = 32'h400e147a; // @[FCLayer.scala 20:24]
  assign mul_8_io_in_a_14 = 32'h40933333; // @[FCLayer.scala 20:24]
  assign mul_8_io_in_a_15 = 32'h3f8a3d70; // @[FCLayer.scala 20:24]
  assign mul_8_io_in_b_0 = io_matB_0; // @[FCLayer.scala 21:24]
  assign mul_8_io_in_b_1 = io_matB_1; // @[FCLayer.scala 21:24]
  assign mul_8_io_in_b_2 = io_matB_2; // @[FCLayer.scala 21:24]
  assign mul_8_io_in_b_3 = io_matB_3; // @[FCLayer.scala 21:24]
  assign mul_8_io_in_b_4 = io_matB_4; // @[FCLayer.scala 21:24]
  assign mul_8_io_in_b_5 = io_matB_5; // @[FCLayer.scala 21:24]
  assign mul_8_io_in_b_6 = io_matB_6; // @[FCLayer.scala 21:24]
  assign mul_8_io_in_b_7 = io_matB_7; // @[FCLayer.scala 21:24]
  assign mul_8_io_in_b_8 = io_matB_8; // @[FCLayer.scala 21:24]
  assign mul_8_io_in_b_9 = io_matB_9; // @[FCLayer.scala 21:24]
  assign mul_8_io_in_b_10 = io_matB_10; // @[FCLayer.scala 21:24]
  assign mul_8_io_in_b_11 = io_matB_11; // @[FCLayer.scala 21:24]
  assign mul_8_io_in_b_12 = io_matB_12; // @[FCLayer.scala 21:24]
  assign mul_8_io_in_b_13 = io_matB_13; // @[FCLayer.scala 21:24]
  assign mul_8_io_in_b_14 = io_matB_14; // @[FCLayer.scala 21:24]
  assign mul_8_io_in_b_15 = io_matB_15; // @[FCLayer.scala 21:24]
  assign fp_adder_8_io_in_a = mul_8_io_out_s; // @[FCLayer.scala 24:24]
  assign fp_adder_8_io_in_b = 32'h40066666; // @[FCLayer.scala 25:24]
  assign mul_9_io_in_a_0 = 32'h4015c28f; // @[FCLayer.scala 20:24]
  assign mul_9_io_in_a_1 = 32'h4007ae14; // @[FCLayer.scala 20:24]
  assign mul_9_io_in_a_2 = 32'h40f47ae1; // @[FCLayer.scala 20:24]
  assign mul_9_io_in_a_3 = 32'h4110a3d7; // @[FCLayer.scala 20:24]
  assign mul_9_io_in_a_4 = 32'h4015c28f; // @[FCLayer.scala 20:24]
  assign mul_9_io_in_a_5 = 32'h3f9d70a3; // @[FCLayer.scala 20:24]
  assign mul_9_io_in_a_6 = 32'h3f9d70a3; // @[FCLayer.scala 20:24]
  assign mul_9_io_in_a_7 = 32'h4087ae14; // @[FCLayer.scala 20:24]
  assign mul_9_io_in_a_8 = 32'h40d1eb85; // @[FCLayer.scala 20:24]
  assign mul_9_io_in_a_9 = 32'h40000000; // @[FCLayer.scala 20:24]
  assign mul_9_io_in_a_10 = 32'h3f800000; // @[FCLayer.scala 20:24]
  assign mul_9_io_in_a_11 = 32'h40400000; // @[FCLayer.scala 20:24]
  assign mul_9_io_in_a_12 = 32'h40800000; // @[FCLayer.scala 20:24]
  assign mul_9_io_in_a_13 = 32'h40a00000; // @[FCLayer.scala 20:24]
  assign mul_9_io_in_a_14 = 32'h40c00000; // @[FCLayer.scala 20:24]
  assign mul_9_io_in_a_15 = 32'h40e00000; // @[FCLayer.scala 20:24]
  assign mul_9_io_in_b_0 = io_matB_0; // @[FCLayer.scala 21:24]
  assign mul_9_io_in_b_1 = io_matB_1; // @[FCLayer.scala 21:24]
  assign mul_9_io_in_b_2 = io_matB_2; // @[FCLayer.scala 21:24]
  assign mul_9_io_in_b_3 = io_matB_3; // @[FCLayer.scala 21:24]
  assign mul_9_io_in_b_4 = io_matB_4; // @[FCLayer.scala 21:24]
  assign mul_9_io_in_b_5 = io_matB_5; // @[FCLayer.scala 21:24]
  assign mul_9_io_in_b_6 = io_matB_6; // @[FCLayer.scala 21:24]
  assign mul_9_io_in_b_7 = io_matB_7; // @[FCLayer.scala 21:24]
  assign mul_9_io_in_b_8 = io_matB_8; // @[FCLayer.scala 21:24]
  assign mul_9_io_in_b_9 = io_matB_9; // @[FCLayer.scala 21:24]
  assign mul_9_io_in_b_10 = io_matB_10; // @[FCLayer.scala 21:24]
  assign mul_9_io_in_b_11 = io_matB_11; // @[FCLayer.scala 21:24]
  assign mul_9_io_in_b_12 = io_matB_12; // @[FCLayer.scala 21:24]
  assign mul_9_io_in_b_13 = io_matB_13; // @[FCLayer.scala 21:24]
  assign mul_9_io_in_b_14 = io_matB_14; // @[FCLayer.scala 21:24]
  assign mul_9_io_in_b_15 = io_matB_15; // @[FCLayer.scala 21:24]
  assign fp_adder_9_io_in_a = mul_9_io_out_s; // @[FCLayer.scala 24:24]
  assign fp_adder_9_io_in_b = 32'h3f800000; // @[FCLayer.scala 25:24]
endmodule
module DigitPrediction(
  input  [31:0] io_input_0,
  input  [31:0] io_input_1,
  input  [31:0] io_input_2,
  input  [31:0] io_input_3,
  input  [31:0] io_input_4,
  input  [31:0] io_input_5,
  input  [31:0] io_input_6,
  input  [31:0] io_input_7,
  input  [31:0] io_input_8,
  input  [31:0] io_input_9,
  output [31:0] io_Digit
);
  wire [31:0] fp1_io_in_a; // @[SoftMax.scala 27:21]
  wire [31:0] fp1_io_in_b; // @[SoftMax.scala 27:21]
  wire [31:0] fp1_io_out_s; // @[SoftMax.scala 27:21]
  wire [31:0] fp2_io_in_a; // @[SoftMax.scala 32:21]
  wire [31:0] fp2_io_in_b; // @[SoftMax.scala 32:21]
  wire [31:0] fp2_io_out_s; // @[SoftMax.scala 32:21]
  wire [31:0] fp3_io_in_a; // @[SoftMax.scala 37:21]
  wire [31:0] fp3_io_in_b; // @[SoftMax.scala 37:21]
  wire [31:0] fp3_io_out_s; // @[SoftMax.scala 37:21]
  wire [31:0] fp4_io_in_a; // @[SoftMax.scala 42:21]
  wire [31:0] fp4_io_in_b; // @[SoftMax.scala 42:21]
  wire [31:0] fp4_io_out_s; // @[SoftMax.scala 42:21]
  wire [31:0] fp5_io_in_a; // @[SoftMax.scala 47:21]
  wire [31:0] fp5_io_in_b; // @[SoftMax.scala 47:21]
  wire [31:0] fp5_io_out_s; // @[SoftMax.scala 47:21]
  wire [31:0] fp6_io_in_a; // @[SoftMax.scala 52:21]
  wire [31:0] fp6_io_in_b; // @[SoftMax.scala 52:21]
  wire [31:0] fp6_io_out_s; // @[SoftMax.scala 52:21]
  wire [31:0] fp7_io_in_a; // @[SoftMax.scala 57:21]
  wire [31:0] fp7_io_in_b; // @[SoftMax.scala 57:21]
  wire [31:0] fp7_io_out_s; // @[SoftMax.scala 57:21]
  wire [31:0] fp8_io_in_a; // @[SoftMax.scala 62:21]
  wire [31:0] fp8_io_in_b; // @[SoftMax.scala 62:21]
  wire [31:0] fp8_io_out_s; // @[SoftMax.scala 62:21]
  wire [31:0] fp9_io_in_a; // @[SoftMax.scala 67:21]
  wire [31:0] fp9_io_in_b; // @[SoftMax.scala 67:21]
  wire [31:0] fp9_io_out_s; // @[SoftMax.scala 67:21]
  wire [31:0] maximum = fp9_io_out_s; // @[SoftMax.scala 22:23 70:13]
  wire [3:0] _GEN_0 = maximum == io_input_8 ? 4'h8 : 4'h9; // @[SoftMax.scala 92:44 93:18 95:18]
  wire [3:0] _GEN_1 = maximum == io_input_7 ? 4'h7 : _GEN_0; // @[SoftMax.scala 90:44 91:18]
  wire [3:0] _GEN_2 = maximum == io_input_6 ? 4'h6 : _GEN_1; // @[SoftMax.scala 88:44 89:18]
  wire [3:0] _GEN_3 = maximum == io_input_5 ? 4'h5 : _GEN_2; // @[SoftMax.scala 86:44 87:18]
  wire [3:0] _GEN_4 = maximum == io_input_4 ? 4'h4 : _GEN_3; // @[SoftMax.scala 84:44 85:18]
  wire [3:0] _GEN_5 = maximum == io_input_3 ? 4'h3 : _GEN_4; // @[SoftMax.scala 82:44 83:18]
  wire [3:0] _GEN_6 = maximum == io_input_2 ? 4'h2 : _GEN_5; // @[SoftMax.scala 80:44 81:18]
  wire [3:0] _GEN_7 = maximum == io_input_1 ? 4'h1 : _GEN_6; // @[SoftMax.scala 78:44 79:18]
  wire [3:0] position = maximum == io_input_0 ? 4'h0 : _GEN_7; // @[SoftMax.scala 76:36 77:18]
  FP_Comparitor fp1 ( // @[SoftMax.scala 27:21]
    .io_in_a(fp1_io_in_a),
    .io_in_b(fp1_io_in_b),
    .io_out_s(fp1_io_out_s)
  );
  FP_Comparitor fp2 ( // @[SoftMax.scala 32:21]
    .io_in_a(fp2_io_in_a),
    .io_in_b(fp2_io_in_b),
    .io_out_s(fp2_io_out_s)
  );
  FP_Comparitor fp3 ( // @[SoftMax.scala 37:21]
    .io_in_a(fp3_io_in_a),
    .io_in_b(fp3_io_in_b),
    .io_out_s(fp3_io_out_s)
  );
  FP_Comparitor fp4 ( // @[SoftMax.scala 42:21]
    .io_in_a(fp4_io_in_a),
    .io_in_b(fp4_io_in_b),
    .io_out_s(fp4_io_out_s)
  );
  FP_Comparitor fp5 ( // @[SoftMax.scala 47:21]
    .io_in_a(fp5_io_in_a),
    .io_in_b(fp5_io_in_b),
    .io_out_s(fp5_io_out_s)
  );
  FP_Comparitor fp6 ( // @[SoftMax.scala 52:21]
    .io_in_a(fp6_io_in_a),
    .io_in_b(fp6_io_in_b),
    .io_out_s(fp6_io_out_s)
  );
  FP_Comparitor fp7 ( // @[SoftMax.scala 57:21]
    .io_in_a(fp7_io_in_a),
    .io_in_b(fp7_io_in_b),
    .io_out_s(fp7_io_out_s)
  );
  FP_Comparitor fp8 ( // @[SoftMax.scala 62:21]
    .io_in_a(fp8_io_in_a),
    .io_in_b(fp8_io_in_b),
    .io_out_s(fp8_io_out_s)
  );
  FP_Comparitor fp9 ( // @[SoftMax.scala 67:21]
    .io_in_a(fp9_io_in_a),
    .io_in_b(fp9_io_in_b),
    .io_out_s(fp9_io_out_s)
  );
  assign io_Digit = {{28'd0}, position}; // @[SoftMax.scala 98:14]
  assign fp1_io_in_a = io_input_0; // @[SoftMax.scala 28:17]
  assign fp1_io_in_b = io_input_1; // @[SoftMax.scala 29:17]
  assign fp2_io_in_a = io_input_2; // @[SoftMax.scala 33:17]
  assign fp2_io_in_b = io_input_3; // @[SoftMax.scala 34:17]
  assign fp3_io_in_a = io_input_4; // @[SoftMax.scala 38:17]
  assign fp3_io_in_b = io_input_5; // @[SoftMax.scala 39:17]
  assign fp4_io_in_a = io_input_6; // @[SoftMax.scala 43:17]
  assign fp4_io_in_b = io_input_7; // @[SoftMax.scala 44:17]
  assign fp5_io_in_a = io_input_8; // @[SoftMax.scala 48:17]
  assign fp5_io_in_b = io_input_9; // @[SoftMax.scala 49:17]
  assign fp6_io_in_a = fp1_io_out_s; // @[SoftMax.scala 14:20 30:10]
  assign fp6_io_in_b = fp2_io_out_s; // @[SoftMax.scala 15:20 35:10]
  assign fp7_io_in_a = fp3_io_out_s; // @[SoftMax.scala 16:20 40:10]
  assign fp7_io_in_b = fp4_io_out_s; // @[SoftMax.scala 17:20 45:10]
  assign fp8_io_in_a = fp6_io_out_s; // @[SoftMax.scala 19:20 55:10]
  assign fp8_io_in_b = fp7_io_out_s; // @[SoftMax.scala 20:20 60:10]
  assign fp9_io_in_a = fp8_io_out_s; // @[SoftMax.scala 21:20 65:10]
  assign fp9_io_in_b = fp5_io_out_s; // @[SoftMax.scala 18:20 50:10]
endmodule
module CNNEngine(
  input         clock,
  input         reset,
  output [31:0] io_Digit
);
  wire [31:0] MatController_io_single_out_0; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_1; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_2; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_3; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_4; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_5; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_6; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_7; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_8; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_9; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_10; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_11; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_12; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_13; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_14; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_15; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_16; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_17; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_18; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_19; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_20; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_21; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_22; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_23; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_24; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_25; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_26; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_27; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_28; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_29; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_30; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_31; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_32; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_33; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_34; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_35; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_36; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_37; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_38; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_39; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_40; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_41; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_42; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_43; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_44; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_45; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_46; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_47; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_48; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_49; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_50; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_51; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_52; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_53; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_54; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_55; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_56; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_57; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_58; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_59; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_60; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_61; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_62; // @[NeuralNetwork.scala 22:31]
  wire [31:0] MatController_io_single_out_63; // @[NeuralNetwork.scala 22:31]
  wire  PoolingControl_clock; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_0; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_1; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_2; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_3; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_4; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_5; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_6; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_7; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_8; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_9; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_10; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_11; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_12; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_13; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_14; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_15; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_16; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_17; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_18; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_19; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_20; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_21; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_22; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_23; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_24; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_25; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_26; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_27; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_28; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_29; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_30; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_31; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_32; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_33; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_34; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_35; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_36; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_37; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_38; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_39; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_40; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_41; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_42; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_43; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_44; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_45; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_46; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_47; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_48; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_49; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_50; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_51; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_52; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_53; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_54; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_55; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_56; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_57; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_58; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_59; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_60; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_61; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_62; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_InputMatrix_63; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_single_out_0; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_single_out_1; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_single_out_2; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_single_out_3; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_single_out_4; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_single_out_5; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_single_out_6; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_single_out_7; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_single_out_8; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_single_out_9; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_single_out_10; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_single_out_11; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_single_out_12; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_single_out_13; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_single_out_14; // @[NeuralNetwork.scala 32:32]
  wire [31:0] PoolingControl_io_single_out_15; // @[NeuralNetwork.scala 32:32]
  wire [31:0] FullyConnected_io_matB_0; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_matB_1; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_matB_2; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_matB_3; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_matB_4; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_matB_5; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_matB_6; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_matB_7; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_matB_8; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_matB_9; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_matB_10; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_matB_11; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_matB_12; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_matB_13; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_matB_14; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_matB_15; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_fC_out_0; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_fC_out_1; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_fC_out_2; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_fC_out_3; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_fC_out_4; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_fC_out_5; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_fC_out_6; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_fC_out_7; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_fC_out_8; // @[NeuralNetwork.scala 39:32]
  wire [31:0] FullyConnected_io_fC_out_9; // @[NeuralNetwork.scala 39:32]
  wire [31:0] SoftMaxModule_io_input_0; // @[NeuralNetwork.scala 55:31]
  wire [31:0] SoftMaxModule_io_input_1; // @[NeuralNetwork.scala 55:31]
  wire [31:0] SoftMaxModule_io_input_2; // @[NeuralNetwork.scala 55:31]
  wire [31:0] SoftMaxModule_io_input_3; // @[NeuralNetwork.scala 55:31]
  wire [31:0] SoftMaxModule_io_input_4; // @[NeuralNetwork.scala 55:31]
  wire [31:0] SoftMaxModule_io_input_5; // @[NeuralNetwork.scala 55:31]
  wire [31:0] SoftMaxModule_io_input_6; // @[NeuralNetwork.scala 55:31]
  wire [31:0] SoftMaxModule_io_input_7; // @[NeuralNetwork.scala 55:31]
  wire [31:0] SoftMaxModule_io_input_8; // @[NeuralNetwork.scala 55:31]
  wire [31:0] SoftMaxModule_io_input_9; // @[NeuralNetwork.scala 55:31]
  wire [31:0] SoftMaxModule_io_Digit; // @[NeuralNetwork.scala 55:31]
  Matrix_Controller MatController ( // @[NeuralNetwork.scala 22:31]
    .io_single_out_0(MatController_io_single_out_0),
    .io_single_out_1(MatController_io_single_out_1),
    .io_single_out_2(MatController_io_single_out_2),
    .io_single_out_3(MatController_io_single_out_3),
    .io_single_out_4(MatController_io_single_out_4),
    .io_single_out_5(MatController_io_single_out_5),
    .io_single_out_6(MatController_io_single_out_6),
    .io_single_out_7(MatController_io_single_out_7),
    .io_single_out_8(MatController_io_single_out_8),
    .io_single_out_9(MatController_io_single_out_9),
    .io_single_out_10(MatController_io_single_out_10),
    .io_single_out_11(MatController_io_single_out_11),
    .io_single_out_12(MatController_io_single_out_12),
    .io_single_out_13(MatController_io_single_out_13),
    .io_single_out_14(MatController_io_single_out_14),
    .io_single_out_15(MatController_io_single_out_15),
    .io_single_out_16(MatController_io_single_out_16),
    .io_single_out_17(MatController_io_single_out_17),
    .io_single_out_18(MatController_io_single_out_18),
    .io_single_out_19(MatController_io_single_out_19),
    .io_single_out_20(MatController_io_single_out_20),
    .io_single_out_21(MatController_io_single_out_21),
    .io_single_out_22(MatController_io_single_out_22),
    .io_single_out_23(MatController_io_single_out_23),
    .io_single_out_24(MatController_io_single_out_24),
    .io_single_out_25(MatController_io_single_out_25),
    .io_single_out_26(MatController_io_single_out_26),
    .io_single_out_27(MatController_io_single_out_27),
    .io_single_out_28(MatController_io_single_out_28),
    .io_single_out_29(MatController_io_single_out_29),
    .io_single_out_30(MatController_io_single_out_30),
    .io_single_out_31(MatController_io_single_out_31),
    .io_single_out_32(MatController_io_single_out_32),
    .io_single_out_33(MatController_io_single_out_33),
    .io_single_out_34(MatController_io_single_out_34),
    .io_single_out_35(MatController_io_single_out_35),
    .io_single_out_36(MatController_io_single_out_36),
    .io_single_out_37(MatController_io_single_out_37),
    .io_single_out_38(MatController_io_single_out_38),
    .io_single_out_39(MatController_io_single_out_39),
    .io_single_out_40(MatController_io_single_out_40),
    .io_single_out_41(MatController_io_single_out_41),
    .io_single_out_42(MatController_io_single_out_42),
    .io_single_out_43(MatController_io_single_out_43),
    .io_single_out_44(MatController_io_single_out_44),
    .io_single_out_45(MatController_io_single_out_45),
    .io_single_out_46(MatController_io_single_out_46),
    .io_single_out_47(MatController_io_single_out_47),
    .io_single_out_48(MatController_io_single_out_48),
    .io_single_out_49(MatController_io_single_out_49),
    .io_single_out_50(MatController_io_single_out_50),
    .io_single_out_51(MatController_io_single_out_51),
    .io_single_out_52(MatController_io_single_out_52),
    .io_single_out_53(MatController_io_single_out_53),
    .io_single_out_54(MatController_io_single_out_54),
    .io_single_out_55(MatController_io_single_out_55),
    .io_single_out_56(MatController_io_single_out_56),
    .io_single_out_57(MatController_io_single_out_57),
    .io_single_out_58(MatController_io_single_out_58),
    .io_single_out_59(MatController_io_single_out_59),
    .io_single_out_60(MatController_io_single_out_60),
    .io_single_out_61(MatController_io_single_out_61),
    .io_single_out_62(MatController_io_single_out_62),
    .io_single_out_63(MatController_io_single_out_63)
  );
  Pooling_Controller PoolingControl ( // @[NeuralNetwork.scala 32:32]
    .clock(PoolingControl_clock),
    .io_InputMatrix_0(PoolingControl_io_InputMatrix_0),
    .io_InputMatrix_1(PoolingControl_io_InputMatrix_1),
    .io_InputMatrix_2(PoolingControl_io_InputMatrix_2),
    .io_InputMatrix_3(PoolingControl_io_InputMatrix_3),
    .io_InputMatrix_4(PoolingControl_io_InputMatrix_4),
    .io_InputMatrix_5(PoolingControl_io_InputMatrix_5),
    .io_InputMatrix_6(PoolingControl_io_InputMatrix_6),
    .io_InputMatrix_7(PoolingControl_io_InputMatrix_7),
    .io_InputMatrix_8(PoolingControl_io_InputMatrix_8),
    .io_InputMatrix_9(PoolingControl_io_InputMatrix_9),
    .io_InputMatrix_10(PoolingControl_io_InputMatrix_10),
    .io_InputMatrix_11(PoolingControl_io_InputMatrix_11),
    .io_InputMatrix_12(PoolingControl_io_InputMatrix_12),
    .io_InputMatrix_13(PoolingControl_io_InputMatrix_13),
    .io_InputMatrix_14(PoolingControl_io_InputMatrix_14),
    .io_InputMatrix_15(PoolingControl_io_InputMatrix_15),
    .io_InputMatrix_16(PoolingControl_io_InputMatrix_16),
    .io_InputMatrix_17(PoolingControl_io_InputMatrix_17),
    .io_InputMatrix_18(PoolingControl_io_InputMatrix_18),
    .io_InputMatrix_19(PoolingControl_io_InputMatrix_19),
    .io_InputMatrix_20(PoolingControl_io_InputMatrix_20),
    .io_InputMatrix_21(PoolingControl_io_InputMatrix_21),
    .io_InputMatrix_22(PoolingControl_io_InputMatrix_22),
    .io_InputMatrix_23(PoolingControl_io_InputMatrix_23),
    .io_InputMatrix_24(PoolingControl_io_InputMatrix_24),
    .io_InputMatrix_25(PoolingControl_io_InputMatrix_25),
    .io_InputMatrix_26(PoolingControl_io_InputMatrix_26),
    .io_InputMatrix_27(PoolingControl_io_InputMatrix_27),
    .io_InputMatrix_28(PoolingControl_io_InputMatrix_28),
    .io_InputMatrix_29(PoolingControl_io_InputMatrix_29),
    .io_InputMatrix_30(PoolingControl_io_InputMatrix_30),
    .io_InputMatrix_31(PoolingControl_io_InputMatrix_31),
    .io_InputMatrix_32(PoolingControl_io_InputMatrix_32),
    .io_InputMatrix_33(PoolingControl_io_InputMatrix_33),
    .io_InputMatrix_34(PoolingControl_io_InputMatrix_34),
    .io_InputMatrix_35(PoolingControl_io_InputMatrix_35),
    .io_InputMatrix_36(PoolingControl_io_InputMatrix_36),
    .io_InputMatrix_37(PoolingControl_io_InputMatrix_37),
    .io_InputMatrix_38(PoolingControl_io_InputMatrix_38),
    .io_InputMatrix_39(PoolingControl_io_InputMatrix_39),
    .io_InputMatrix_40(PoolingControl_io_InputMatrix_40),
    .io_InputMatrix_41(PoolingControl_io_InputMatrix_41),
    .io_InputMatrix_42(PoolingControl_io_InputMatrix_42),
    .io_InputMatrix_43(PoolingControl_io_InputMatrix_43),
    .io_InputMatrix_44(PoolingControl_io_InputMatrix_44),
    .io_InputMatrix_45(PoolingControl_io_InputMatrix_45),
    .io_InputMatrix_46(PoolingControl_io_InputMatrix_46),
    .io_InputMatrix_47(PoolingControl_io_InputMatrix_47),
    .io_InputMatrix_48(PoolingControl_io_InputMatrix_48),
    .io_InputMatrix_49(PoolingControl_io_InputMatrix_49),
    .io_InputMatrix_50(PoolingControl_io_InputMatrix_50),
    .io_InputMatrix_51(PoolingControl_io_InputMatrix_51),
    .io_InputMatrix_52(PoolingControl_io_InputMatrix_52),
    .io_InputMatrix_53(PoolingControl_io_InputMatrix_53),
    .io_InputMatrix_54(PoolingControl_io_InputMatrix_54),
    .io_InputMatrix_55(PoolingControl_io_InputMatrix_55),
    .io_InputMatrix_56(PoolingControl_io_InputMatrix_56),
    .io_InputMatrix_57(PoolingControl_io_InputMatrix_57),
    .io_InputMatrix_58(PoolingControl_io_InputMatrix_58),
    .io_InputMatrix_59(PoolingControl_io_InputMatrix_59),
    .io_InputMatrix_60(PoolingControl_io_InputMatrix_60),
    .io_InputMatrix_61(PoolingControl_io_InputMatrix_61),
    .io_InputMatrix_62(PoolingControl_io_InputMatrix_62),
    .io_InputMatrix_63(PoolingControl_io_InputMatrix_63),
    .io_single_out_0(PoolingControl_io_single_out_0),
    .io_single_out_1(PoolingControl_io_single_out_1),
    .io_single_out_2(PoolingControl_io_single_out_2),
    .io_single_out_3(PoolingControl_io_single_out_3),
    .io_single_out_4(PoolingControl_io_single_out_4),
    .io_single_out_5(PoolingControl_io_single_out_5),
    .io_single_out_6(PoolingControl_io_single_out_6),
    .io_single_out_7(PoolingControl_io_single_out_7),
    .io_single_out_8(PoolingControl_io_single_out_8),
    .io_single_out_9(PoolingControl_io_single_out_9),
    .io_single_out_10(PoolingControl_io_single_out_10),
    .io_single_out_11(PoolingControl_io_single_out_11),
    .io_single_out_12(PoolingControl_io_single_out_12),
    .io_single_out_13(PoolingControl_io_single_out_13),
    .io_single_out_14(PoolingControl_io_single_out_14),
    .io_single_out_15(PoolingControl_io_single_out_15)
  );
  FC FullyConnected ( // @[NeuralNetwork.scala 39:32]
    .io_matB_0(FullyConnected_io_matB_0),
    .io_matB_1(FullyConnected_io_matB_1),
    .io_matB_2(FullyConnected_io_matB_2),
    .io_matB_3(FullyConnected_io_matB_3),
    .io_matB_4(FullyConnected_io_matB_4),
    .io_matB_5(FullyConnected_io_matB_5),
    .io_matB_6(FullyConnected_io_matB_6),
    .io_matB_7(FullyConnected_io_matB_7),
    .io_matB_8(FullyConnected_io_matB_8),
    .io_matB_9(FullyConnected_io_matB_9),
    .io_matB_10(FullyConnected_io_matB_10),
    .io_matB_11(FullyConnected_io_matB_11),
    .io_matB_12(FullyConnected_io_matB_12),
    .io_matB_13(FullyConnected_io_matB_13),
    .io_matB_14(FullyConnected_io_matB_14),
    .io_matB_15(FullyConnected_io_matB_15),
    .io_fC_out_0(FullyConnected_io_fC_out_0),
    .io_fC_out_1(FullyConnected_io_fC_out_1),
    .io_fC_out_2(FullyConnected_io_fC_out_2),
    .io_fC_out_3(FullyConnected_io_fC_out_3),
    .io_fC_out_4(FullyConnected_io_fC_out_4),
    .io_fC_out_5(FullyConnected_io_fC_out_5),
    .io_fC_out_6(FullyConnected_io_fC_out_6),
    .io_fC_out_7(FullyConnected_io_fC_out_7),
    .io_fC_out_8(FullyConnected_io_fC_out_8),
    .io_fC_out_9(FullyConnected_io_fC_out_9)
  );
  DigitPrediction SoftMaxModule ( // @[NeuralNetwork.scala 55:31]
    .io_input_0(SoftMaxModule_io_input_0),
    .io_input_1(SoftMaxModule_io_input_1),
    .io_input_2(SoftMaxModule_io_input_2),
    .io_input_3(SoftMaxModule_io_input_3),
    .io_input_4(SoftMaxModule_io_input_4),
    .io_input_5(SoftMaxModule_io_input_5),
    .io_input_6(SoftMaxModule_io_input_6),
    .io_input_7(SoftMaxModule_io_input_7),
    .io_input_8(SoftMaxModule_io_input_8),
    .io_input_9(SoftMaxModule_io_input_9),
    .io_Digit(SoftMaxModule_io_Digit)
  );
  assign io_Digit = SoftMaxModule_io_Digit; // @[NeuralNetwork.scala 60:14]
  assign PoolingControl_clock = clock;
  assign PoolingControl_io_InputMatrix_0 = MatController_io_single_out_0; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_1 = MatController_io_single_out_1; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_2 = MatController_io_single_out_2; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_3 = MatController_io_single_out_3; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_4 = MatController_io_single_out_4; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_5 = MatController_io_single_out_5; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_6 = MatController_io_single_out_6; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_7 = MatController_io_single_out_7; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_8 = MatController_io_single_out_8; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_9 = MatController_io_single_out_9; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_10 = MatController_io_single_out_10; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_11 = MatController_io_single_out_11; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_12 = MatController_io_single_out_12; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_13 = MatController_io_single_out_13; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_14 = MatController_io_single_out_14; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_15 = MatController_io_single_out_15; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_16 = MatController_io_single_out_16; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_17 = MatController_io_single_out_17; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_18 = MatController_io_single_out_18; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_19 = MatController_io_single_out_19; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_20 = MatController_io_single_out_20; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_21 = MatController_io_single_out_21; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_22 = MatController_io_single_out_22; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_23 = MatController_io_single_out_23; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_24 = MatController_io_single_out_24; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_25 = MatController_io_single_out_25; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_26 = MatController_io_single_out_26; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_27 = MatController_io_single_out_27; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_28 = MatController_io_single_out_28; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_29 = MatController_io_single_out_29; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_30 = MatController_io_single_out_30; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_31 = MatController_io_single_out_31; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_32 = MatController_io_single_out_32; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_33 = MatController_io_single_out_33; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_34 = MatController_io_single_out_34; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_35 = MatController_io_single_out_35; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_36 = MatController_io_single_out_36; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_37 = MatController_io_single_out_37; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_38 = MatController_io_single_out_38; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_39 = MatController_io_single_out_39; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_40 = MatController_io_single_out_40; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_41 = MatController_io_single_out_41; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_42 = MatController_io_single_out_42; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_43 = MatController_io_single_out_43; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_44 = MatController_io_single_out_44; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_45 = MatController_io_single_out_45; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_46 = MatController_io_single_out_46; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_47 = MatController_io_single_out_47; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_48 = MatController_io_single_out_48; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_49 = MatController_io_single_out_49; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_50 = MatController_io_single_out_50; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_51 = MatController_io_single_out_51; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_52 = MatController_io_single_out_52; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_53 = MatController_io_single_out_53; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_54 = MatController_io_single_out_54; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_55 = MatController_io_single_out_55; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_56 = MatController_io_single_out_56; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_57 = MatController_io_single_out_57; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_58 = MatController_io_single_out_58; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_59 = MatController_io_single_out_59; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_60 = MatController_io_single_out_60; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_61 = MatController_io_single_out_61; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_62 = MatController_io_single_out_62; // @[NeuralNetwork.scala 35:40]
  assign PoolingControl_io_InputMatrix_63 = MatController_io_single_out_63; // @[NeuralNetwork.scala 35:40]
  assign FullyConnected_io_matB_0 = PoolingControl_io_single_out_0; // @[NeuralNetwork.scala 42:33]
  assign FullyConnected_io_matB_1 = PoolingControl_io_single_out_1; // @[NeuralNetwork.scala 42:33]
  assign FullyConnected_io_matB_2 = PoolingControl_io_single_out_2; // @[NeuralNetwork.scala 42:33]
  assign FullyConnected_io_matB_3 = PoolingControl_io_single_out_3; // @[NeuralNetwork.scala 42:33]
  assign FullyConnected_io_matB_4 = PoolingControl_io_single_out_4; // @[NeuralNetwork.scala 42:33]
  assign FullyConnected_io_matB_5 = PoolingControl_io_single_out_5; // @[NeuralNetwork.scala 42:33]
  assign FullyConnected_io_matB_6 = PoolingControl_io_single_out_6; // @[NeuralNetwork.scala 42:33]
  assign FullyConnected_io_matB_7 = PoolingControl_io_single_out_7; // @[NeuralNetwork.scala 42:33]
  assign FullyConnected_io_matB_8 = PoolingControl_io_single_out_8; // @[NeuralNetwork.scala 42:33]
  assign FullyConnected_io_matB_9 = PoolingControl_io_single_out_9; // @[NeuralNetwork.scala 42:33]
  assign FullyConnected_io_matB_10 = PoolingControl_io_single_out_10; // @[NeuralNetwork.scala 42:33]
  assign FullyConnected_io_matB_11 = PoolingControl_io_single_out_11; // @[NeuralNetwork.scala 42:33]
  assign FullyConnected_io_matB_12 = PoolingControl_io_single_out_12; // @[NeuralNetwork.scala 42:33]
  assign FullyConnected_io_matB_13 = PoolingControl_io_single_out_13; // @[NeuralNetwork.scala 42:33]
  assign FullyConnected_io_matB_14 = PoolingControl_io_single_out_14; // @[NeuralNetwork.scala 42:33]
  assign FullyConnected_io_matB_15 = PoolingControl_io_single_out_15; // @[NeuralNetwork.scala 42:33]
  assign SoftMaxModule_io_input_0 = FullyConnected_io_fC_out_0; // @[NeuralNetwork.scala 58:33]
  assign SoftMaxModule_io_input_1 = FullyConnected_io_fC_out_1; // @[NeuralNetwork.scala 58:33]
  assign SoftMaxModule_io_input_2 = FullyConnected_io_fC_out_2; // @[NeuralNetwork.scala 58:33]
  assign SoftMaxModule_io_input_3 = FullyConnected_io_fC_out_3; // @[NeuralNetwork.scala 58:33]
  assign SoftMaxModule_io_input_4 = FullyConnected_io_fC_out_4; // @[NeuralNetwork.scala 58:33]
  assign SoftMaxModule_io_input_5 = FullyConnected_io_fC_out_5; // @[NeuralNetwork.scala 58:33]
  assign SoftMaxModule_io_input_6 = FullyConnected_io_fC_out_6; // @[NeuralNetwork.scala 58:33]
  assign SoftMaxModule_io_input_7 = FullyConnected_io_fC_out_7; // @[NeuralNetwork.scala 58:33]
  assign SoftMaxModule_io_input_8 = FullyConnected_io_fC_out_8; // @[NeuralNetwork.scala 58:33]
  assign SoftMaxModule_io_input_9 = FullyConnected_io_fC_out_9; // @[NeuralNetwork.scala 58:33]
endmodule

